                      .MU0_EFPGA_MATHB_COEF_DATA_23_(MU0_EFPGA_MATHB_COEF_DATA[23]),
                      .MU0_EFPGA_MATHB_COEF_DATA_22_(MU0_EFPGA_MATHB_COEF_DATA[22]),
                      .MU0_EFPGA_MATHB_COEF_DATA_13_(MU0_EFPGA_MATHB_COEF_DATA[13]),
                      .MU0_EFPGA_MATHB_COEF_DATA_12_(MU0_EFPGA_MATHB_COEF_DATA[12]),
                      .MU0_EFPGA_MATHB_COEF_DATA_11_(MU0_EFPGA_MATHB_COEF_DATA[11]),
                      .MU0_EFPGA_MATHB_COEF_DATA_10_(MU0_EFPGA_MATHB_COEF_DATA[10]),
                      .MU0_EFPGA_MATHB_COEF_DATA_9_(MU0_EFPGA_MATHB_COEF_DATA[9]),
                      .MU0_EFPGA_MATHB_COEF_DATA_8_(MU0_EFPGA_MATHB_COEF_DATA[8]),
                      .MU0_EFPGA_MATHB_COEF_DATA_7_(MU0_EFPGA_MATHB_COEF_DATA[7]),
                      .MU0_EFPGA_MATHB_COEF_DATA_6_(MU0_EFPGA_MATHB_COEF_DATA[6]),
                      .MU0_EFPGA_MATHB_COEF_DATA_21_(MU0_EFPGA_MATHB_COEF_DATA[21]),
                      .MU0_EFPGA_MATHB_COEF_DATA_20_(MU0_EFPGA_MATHB_COEF_DATA[20]),
                      .MU0_EFPGA_MATHB_COEF_DATA_19_(MU0_EFPGA_MATHB_COEF_DATA[19]),
                      .MU0_EFPGA_MATHB_COEF_DATA_18_(MU0_EFPGA_MATHB_COEF_DATA[18]),
                      .MU0_EFPGA_MATHB_COEF_DATA_17_(MU0_EFPGA_MATHB_COEF_DATA[17]),
                      .MU0_EFPGA_MATHB_COEF_DATA_16_(MU0_EFPGA_MATHB_COEF_DATA[16]),
                      .MU0_EFPGA_MATHB_COEF_DATA_15_(MU0_EFPGA_MATHB_COEF_DATA[15]),
                      .MU0_EFPGA_MATHB_COEF_DATA_14_(MU0_EFPGA_MATHB_COEF_DATA[14]),
                      .MU0_EFPGA_MATHB_COEF_DATA_5_(MU0_EFPGA_MATHB_COEF_DATA[5]),
                      .MU0_EFPGA_MATHB_COEF_DATA_4_(MU0_EFPGA_MATHB_COEF_DATA[4]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_31_(MU0_EFPGA_TPRAM_COEF_W_DATA[31]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_30_(MU0_EFPGA_TPRAM_COEF_W_DATA[30]),
                      .MU0_EFPGA_MATHB_COEF_DATA_3_(MU0_EFPGA_MATHB_COEF_DATA[3]),
                      .MU0_EFPGA_MATHB_COEF_DATA_2_(MU0_EFPGA_MATHB_COEF_DATA[2]),
                      .MU0_EFPGA_MATHB_COEF_DATA_1_(MU0_EFPGA_MATHB_COEF_DATA[1]),
                      .MU0_EFPGA_MATHB_COEF_DATA_0_(MU0_EFPGA_MATHB_COEF_DATA[0]),
                      .MU0_EFPGA_MATHB_DATAOUT_SEL_1_(MU0_EFPGA_MATHB_DATAOUT_SEL[1]),
                      .MU0_EFPGA_MATHB_DATAOUT_SEL_0_(MU0_EFPGA_MATHB_DATAOUT_SEL[0]),
                      .MU0_EFPGA_TPRAM_COEF_W_MODE_1_(MU0_EFPGA_TPRAM_COEF_W_MODE[1]),
                      .MU0_EFPGA_TPRAM_COEF_W_MODE_0_(MU0_EFPGA_TPRAM_COEF_W_MODE[0]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_29_(MU0_EFPGA_TPRAM_COEF_W_DATA[29]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_28_(MU0_EFPGA_TPRAM_COEF_W_DATA[28]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_19_(MU0_EFPGA_TPRAM_COEF_W_DATA[19]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_18_(MU0_EFPGA_TPRAM_COEF_W_DATA[18]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_17_(MU0_EFPGA_TPRAM_COEF_W_DATA[17]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_16_(MU0_EFPGA_TPRAM_COEF_W_DATA[16]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_15_(MU0_EFPGA_TPRAM_COEF_W_DATA[15]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_14_(MU0_EFPGA_TPRAM_COEF_W_DATA[14]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_13_(MU0_EFPGA_TPRAM_COEF_W_DATA[13]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_12_(MU0_EFPGA_TPRAM_COEF_W_DATA[12]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_27_(MU0_EFPGA_TPRAM_COEF_W_DATA[27]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_26_(MU0_EFPGA_TPRAM_COEF_W_DATA[26]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_25_(MU0_EFPGA_TPRAM_COEF_W_DATA[25]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_24_(MU0_EFPGA_TPRAM_COEF_W_DATA[24]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_23_(MU0_EFPGA_TPRAM_COEF_W_DATA[23]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_22_(MU0_EFPGA_TPRAM_COEF_W_DATA[22]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_21_(MU0_EFPGA_TPRAM_COEF_W_DATA[21]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_20_(MU0_EFPGA_TPRAM_COEF_W_DATA[20]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_11_(MU0_EFPGA_TPRAM_COEF_W_DATA[11]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_10_(MU0_EFPGA_TPRAM_COEF_W_DATA[10]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_1_(MU0_EFPGA_TPRAM_COEF_W_DATA[1]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_0_(MU0_EFPGA_TPRAM_COEF_W_DATA[0]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_9_(MU0_EFPGA_TPRAM_COEF_W_DATA[9]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_8_(MU0_EFPGA_TPRAM_COEF_W_DATA[8]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_7_(MU0_EFPGA_TPRAM_COEF_W_DATA[7]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_6_(MU0_EFPGA_TPRAM_COEF_W_DATA[6]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_5_(MU0_EFPGA_TPRAM_COEF_W_DATA[5]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_4_(MU0_EFPGA_TPRAM_COEF_W_DATA[4]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_3_(MU0_EFPGA_TPRAM_COEF_W_DATA[3]),
                      .MU0_EFPGA_TPRAM_COEF_W_DATA_2_(MU0_EFPGA_TPRAM_COEF_W_DATA[2]),
                      .MU0_EFPGA_TPRAM_COEF_W_CLK(MU0_EFPGA_TPRAM_COEF_W_CLK),
                      .MU0_EFPGA_TPRAM_COEF_W_ADDR_11_(MU0_EFPGA_TPRAM_COEF_W_ADDR[11]),
                      .MU0_EFPGA_TPRAM_COEF_W_ADDR_2_(MU0_EFPGA_TPRAM_COEF_W_ADDR[2]),
                      .MU0_EFPGA_TPRAM_COEF_W_ADDR_1_(MU0_EFPGA_TPRAM_COEF_W_ADDR[1]),
                      .MU0_EFPGA_TPRAM_COEF_W_ADDR_0_(MU0_EFPGA_TPRAM_COEF_W_ADDR[0]),
                      .MU0_EFPGA_TPRAM_COEF_WE(MU0_EFPGA_TPRAM_COEF_WE),
                      .MU0_EFPGA_TPRAM_COEF_WDSEL(MU0_EFPGA_TPRAM_COEF_WDSEL),
                      .MU0_EFPGA_TPRAM_COEF_R_MODE_1_(MU0_EFPGA_TPRAM_COEF_R_MODE[1]),
                      .MU0_EFPGA_TPRAM_COEF_R_MODE_0_(MU0_EFPGA_TPRAM_COEF_R_MODE[0]),
                      .MU0_EFPGA_TPRAM_COEF_R_CLK(MU0_EFPGA_TPRAM_COEF_R_CLK),
                      .MU0_EFPGA_TPRAM_COEF_W_ADDR_10_(MU0_EFPGA_TPRAM_COEF_W_ADDR[10]),
                      .MU0_EFPGA_TPRAM_COEF_W_ADDR_9_(MU0_EFPGA_TPRAM_COEF_W_ADDR[9]),
                      .MU0_EFPGA_TPRAM_COEF_W_ADDR_8_(MU0_EFPGA_TPRAM_COEF_W_ADDR[8]),
                      .MU0_EFPGA_TPRAM_COEF_W_ADDR_7_(MU0_EFPGA_TPRAM_COEF_W_ADDR[7]),
                      .MU0_EFPGA_TPRAM_COEF_W_ADDR_6_(MU0_EFPGA_TPRAM_COEF_W_ADDR[6]),
                      .MU0_EFPGA_TPRAM_COEF_W_ADDR_5_(MU0_EFPGA_TPRAM_COEF_W_ADDR[5]),
                      .MU0_EFPGA_TPRAM_COEF_W_ADDR_4_(MU0_EFPGA_TPRAM_COEF_W_ADDR[4]),
                      .MU0_EFPGA_TPRAM_COEF_W_ADDR_3_(MU0_EFPGA_TPRAM_COEF_W_ADDR[3]),
                      .MU0_EFPGA_TPRAM_COEF_R_ADDR_11_(MU0_EFPGA_TPRAM_COEF_R_ADDR[11]),
                      .MU0_EFPGA_TPRAM_COEF_R_ADDR_10_(MU0_EFPGA_TPRAM_COEF_R_ADDR[10]),
                      .MU0_EFPGA_TPRAM_COEF_R_ADDR_1_(MU0_EFPGA_TPRAM_COEF_R_ADDR[1]),
                      .MU0_EFPGA_TPRAM_COEF_R_ADDR_0_(MU0_EFPGA_TPRAM_COEF_R_ADDR[0]),
                      .MU0_EFPGA_TPRAM_COEF_R_ADDR_9_(MU0_EFPGA_TPRAM_COEF_R_ADDR[9]),
                      .MU0_EFPGA_TPRAM_COEF_R_ADDR_8_(MU0_EFPGA_TPRAM_COEF_R_ADDR[8]),
                      .MU0_EFPGA_TPRAM_COEF_R_ADDR_7_(MU0_EFPGA_TPRAM_COEF_R_ADDR[7]),
                      .MU0_EFPGA_TPRAM_COEF_R_ADDR_6_(MU0_EFPGA_TPRAM_COEF_R_ADDR[6]),
                      .MU0_EFPGA_TPRAM_COEF_R_ADDR_5_(MU0_EFPGA_TPRAM_COEF_R_ADDR[5]),
                      .MU0_EFPGA_TPRAM_COEF_R_ADDR_4_(MU0_EFPGA_TPRAM_COEF_R_ADDR[4]),
                      .MU0_EFPGA_TPRAM_COEF_R_ADDR_3_(MU0_EFPGA_TPRAM_COEF_R_ADDR[3]),
                      .MU0_EFPGA_TPRAM_COEF_R_ADDR_2_(MU0_EFPGA_TPRAM_COEF_R_ADDR[2]),
                      .MU0_EFPGA_TPRAM_COEF_POWERDN(MU0_EFPGA_TPRAM_COEF_POWERDN),
                      .MU1_EFPGA_TPRAM_OPER_W_MODE_1_(MU1_EFPGA_TPRAM_OPER_W_MODE[1]),
                      .MU1_EFPGA_TPRAM_OPER_W_MODE_0_(MU1_EFPGA_TPRAM_OPER_W_MODE[0]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_23_(MU1_EFPGA_TPRAM_OPER_W_DATA[23]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_22_(MU1_EFPGA_TPRAM_OPER_W_DATA[22]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_31_(MU1_EFPGA_TPRAM_OPER_W_DATA[31]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_30_(MU1_EFPGA_TPRAM_OPER_W_DATA[30]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_29_(MU1_EFPGA_TPRAM_OPER_W_DATA[29]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_28_(MU1_EFPGA_TPRAM_OPER_W_DATA[28]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_27_(MU1_EFPGA_TPRAM_OPER_W_DATA[27]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_26_(MU1_EFPGA_TPRAM_OPER_W_DATA[26]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_25_(MU1_EFPGA_TPRAM_OPER_W_DATA[25]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_24_(MU1_EFPGA_TPRAM_OPER_W_DATA[24]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_21_(MU1_EFPGA_TPRAM_OPER_W_DATA[21]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_20_(MU1_EFPGA_TPRAM_OPER_W_DATA[20]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_11_(MU1_EFPGA_TPRAM_OPER_W_DATA[11]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_10_(MU1_EFPGA_TPRAM_OPER_W_DATA[10]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_9_(MU1_EFPGA_TPRAM_OPER_W_DATA[9]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_8_(MU1_EFPGA_TPRAM_OPER_W_DATA[8]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_7_(MU1_EFPGA_TPRAM_OPER_W_DATA[7]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_6_(MU1_EFPGA_TPRAM_OPER_W_DATA[6]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_5_(MU1_EFPGA_TPRAM_OPER_W_DATA[5]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_4_(MU1_EFPGA_TPRAM_OPER_W_DATA[4]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_19_(MU1_EFPGA_TPRAM_OPER_W_DATA[19]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_18_(MU1_EFPGA_TPRAM_OPER_W_DATA[18]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_17_(MU1_EFPGA_TPRAM_OPER_W_DATA[17]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_16_(MU1_EFPGA_TPRAM_OPER_W_DATA[16]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_15_(MU1_EFPGA_TPRAM_OPER_W_DATA[15]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_14_(MU1_EFPGA_TPRAM_OPER_W_DATA[14]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_13_(MU1_EFPGA_TPRAM_OPER_W_DATA[13]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_12_(MU1_EFPGA_TPRAM_OPER_W_DATA[12]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_3_(MU1_EFPGA_TPRAM_OPER_W_DATA[3]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_2_(MU1_EFPGA_TPRAM_OPER_W_DATA[2]),
                      .MU1_EFPGA_TPRAM_OPER_W_ADDR_6_(MU1_EFPGA_TPRAM_OPER_W_ADDR[6]),
                      .MU1_EFPGA_TPRAM_OPER_W_ADDR_5_(MU1_EFPGA_TPRAM_OPER_W_ADDR[5]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_1_(MU1_EFPGA_TPRAM_OPER_W_DATA[1]),
                      .MU1_EFPGA_TPRAM_OPER_W_DATA_0_(MU1_EFPGA_TPRAM_OPER_W_DATA[0]),
                      .MU1_EFPGA_TPRAM_OPER_W_CLK(MU1_EFPGA_TPRAM_OPER_W_CLK),
                      .MU1_EFPGA_TPRAM_OPER_W_ADDR_11_(MU1_EFPGA_TPRAM_OPER_W_ADDR[11]),
                      .MU1_EFPGA_TPRAM_OPER_W_ADDR_10_(MU1_EFPGA_TPRAM_OPER_W_ADDR[10]),
                      .MU1_EFPGA_TPRAM_OPER_W_ADDR_9_(MU1_EFPGA_TPRAM_OPER_W_ADDR[9]),
                      .MU1_EFPGA_TPRAM_OPER_W_ADDR_8_(MU1_EFPGA_TPRAM_OPER_W_ADDR[8]),
                      .MU1_EFPGA_TPRAM_OPER_W_ADDR_7_(MU1_EFPGA_TPRAM_OPER_W_ADDR[7]),
                      .MU1_EFPGA_TPRAM_OPER_W_ADDR_4_(MU1_EFPGA_TPRAM_OPER_W_ADDR[4]),
                      .MU1_EFPGA_TPRAM_OPER_W_ADDR_3_(MU1_EFPGA_TPRAM_OPER_W_ADDR[3]),
                      .MU1_EFPGA_TPRAM_OPER_R_ADDR_11_(MU1_EFPGA_TPRAM_OPER_R_ADDR[11]),
                      .MU1_EFPGA_TPRAM_OPER_R_ADDR_10_(MU1_EFPGA_TPRAM_OPER_R_ADDR[10]),
                      .MU1_EFPGA_TPRAM_OPER_R_ADDR_9_(MU1_EFPGA_TPRAM_OPER_R_ADDR[9]),
                      .MU1_EFPGA_TPRAM_OPER_R_ADDR_8_(MU1_EFPGA_TPRAM_OPER_R_ADDR[8]),
                      .MU1_EFPGA_TPRAM_OPER_R_ADDR_7_(MU1_EFPGA_TPRAM_OPER_R_ADDR[7]),
                      .MU1_EFPGA_TPRAM_OPER_R_ADDR_6_(MU1_EFPGA_TPRAM_OPER_R_ADDR[6]),
                      .MU1_EFPGA_TPRAM_OPER_R_ADDR_5_(MU1_EFPGA_TPRAM_OPER_R_ADDR[5]),
                      .MU1_EFPGA_TPRAM_OPER_R_ADDR_4_(MU1_EFPGA_TPRAM_OPER_R_ADDR[4]),
                      .MU1_EFPGA_TPRAM_OPER_W_ADDR_2_(MU1_EFPGA_TPRAM_OPER_W_ADDR[2]),
                      .MU1_EFPGA_TPRAM_OPER_W_ADDR_1_(MU1_EFPGA_TPRAM_OPER_W_ADDR[1]),
                      .MU1_EFPGA_TPRAM_OPER_W_ADDR_0_(MU1_EFPGA_TPRAM_OPER_W_ADDR[0]),
                      .MU1_EFPGA_TPRAM_OPER_WE(MU1_EFPGA_TPRAM_OPER_WE),
                      .MU1_EFPGA_TPRAM_OPER_WDSEL(MU1_EFPGA_TPRAM_OPER_WDSEL),
                      .MU1_EFPGA_TPRAM_OPER_R_MODE_1_(MU1_EFPGA_TPRAM_OPER_R_MODE[1]),
                      .MU1_EFPGA_TPRAM_OPER_R_MODE_0_(MU1_EFPGA_TPRAM_OPER_R_MODE[0]),
                      .MU1_EFPGA_TPRAM_OPER_R_CLK(MU1_EFPGA_TPRAM_OPER_R_CLK),
                      .MU1_EFPGA_TPRAM_OPER_R_ADDR_3_(MU1_EFPGA_TPRAM_OPER_R_ADDR[3]),
                      .MU1_EFPGA_TPRAM_OPER_R_ADDR_2_(MU1_EFPGA_TPRAM_OPER_R_ADDR[2]),
                      .MU1_EFPGA_MATHB_MAC_OUT_SEL_2_(MU1_EFPGA_MATHB_MAC_OUT_SEL[2]),
                      .MU1_EFPGA_MATHB_MAC_OUT_SEL_1_(MU1_EFPGA_MATHB_MAC_OUT_SEL[1]),
                      .MU1_EFPGA_TPRAM_OPER_R_ADDR_1_(MU1_EFPGA_TPRAM_OPER_R_ADDR[1]),
                      .MU1_EFPGA_TPRAM_OPER_R_ADDR_0_(MU1_EFPGA_TPRAM_OPER_R_ADDR[0]),
                      .MU1_EFPGA_TPRAM_OPER_POWERDN(MU1_EFPGA_TPRAM_OPER_POWERDN),
                      .MU1_EFPGA2MATHB_CLK(MU1_EFPGA2MATHB_CLK),
                      .MU1_EFPGA_MATHB_CLK_EN(MU1_EFPGA_MATHB_CLK_EN),
                      .MU1_EFPGA_MATHB_MAC_OUT_SEL_5_(MU1_EFPGA_MATHB_MAC_OUT_SEL[5]),
                      .MU1_EFPGA_MATHB_MAC_OUT_SEL_4_(MU1_EFPGA_MATHB_MAC_OUT_SEL[4]),
                      .MU1_EFPGA_MATHB_MAC_OUT_SEL_3_(MU1_EFPGA_MATHB_MAC_OUT_SEL[3]),
                      .MU1_EFPGA_MATHB_MAC_OUT_SEL_0_(MU1_EFPGA_MATHB_MAC_OUT_SEL[0]),
                      .MU1_EFPGA_MATHB_MAC_ACC_SAT(MU1_EFPGA_MATHB_MAC_ACC_SAT),
                      .MU1_EFPGA_MATHB_OPER_DATA_26_(MU1_EFPGA_MATHB_OPER_DATA[26]),
                      .MU1_EFPGA_MATHB_OPER_DATA_25_(MU1_EFPGA_MATHB_OPER_DATA[25]),
                      .MU1_EFPGA_MATHB_OPER_DATA_24_(MU1_EFPGA_MATHB_OPER_DATA[24]),
                      .MU1_EFPGA_MATHB_OPER_DATA_23_(MU1_EFPGA_MATHB_OPER_DATA[23]),
                      .MU1_EFPGA_MATHB_OPER_DATA_22_(MU1_EFPGA_MATHB_OPER_DATA[22]),
                      .MU1_EFPGA_MATHB_OPER_DATA_21_(MU1_EFPGA_MATHB_OPER_DATA[21]),
                      .MU1_EFPGA_MATHB_OPER_DATA_20_(MU1_EFPGA_MATHB_OPER_DATA[20]),
                      .MU1_EFPGA_MATHB_OPER_DATA_19_(MU1_EFPGA_MATHB_OPER_DATA[19]),
                      .MU1_EFPGA_MATHB_MAC_ACC_RND(MU1_EFPGA_MATHB_MAC_ACC_RND),
                      .MU1_EFPGA_MATHB_MAC_ACC_CLEAR(MU1_EFPGA_MATHB_MAC_ACC_CLEAR),
                      .MU1_EFPGA_MATHB_OPER_SEL(MU1_EFPGA_MATHB_OPER_SEL),
                      .MU1_EFPGA_MATHB_OPER_DATA_31_(MU1_EFPGA_MATHB_OPER_DATA[31]),
                      .MU1_EFPGA_MATHB_OPER_DATA_30_(MU1_EFPGA_MATHB_OPER_DATA[30]),
                      .MU1_EFPGA_MATHB_OPER_DATA_29_(MU1_EFPGA_MATHB_OPER_DATA[29]),
                      .MU1_EFPGA_MATHB_OPER_DATA_28_(MU1_EFPGA_MATHB_OPER_DATA[28]),
                      .MU1_EFPGA_MATHB_OPER_DATA_27_(MU1_EFPGA_MATHB_OPER_DATA[27]),
                      .MU1_EFPGA_MATHB_OPER_DATA_18_(MU1_EFPGA_MATHB_OPER_DATA[18]),
                      .MU1_EFPGA_MATHB_OPER_DATA_17_(MU1_EFPGA_MATHB_OPER_DATA[17]),
                      .MU1_EFPGA_MATHB_OPER_DATA_8_(MU1_EFPGA_MATHB_OPER_DATA[8]),
                      .MU1_EFPGA_MATHB_OPER_DATA_7_(MU1_EFPGA_MATHB_OPER_DATA[7]),
                      .MU1_EFPGA_MATHB_OPER_DATA_16_(MU1_EFPGA_MATHB_OPER_DATA[16]),
                      .MU1_EFPGA_MATHB_OPER_DATA_15_(MU1_EFPGA_MATHB_OPER_DATA[15]),
                      .MU1_EFPGA_MATHB_OPER_DATA_14_(MU1_EFPGA_MATHB_OPER_DATA[14]),
                      .MU1_EFPGA_MATHB_OPER_DATA_13_(MU1_EFPGA_MATHB_OPER_DATA[13]),
                      .MU1_EFPGA_MATHB_OPER_DATA_12_(MU1_EFPGA_MATHB_OPER_DATA[12]),
                      .MU1_EFPGA_MATHB_OPER_DATA_11_(MU1_EFPGA_MATHB_OPER_DATA[11]),
                      .MU1_EFPGA_MATHB_OPER_DATA_10_(MU1_EFPGA_MATHB_OPER_DATA[10]),
                      .MU1_EFPGA_MATHB_OPER_DATA_9_(MU1_EFPGA_MATHB_OPER_DATA[9]),
                      .MU1_EFPGA_MATHB_OPER_DATA_6_(MU1_EFPGA_MATHB_OPER_DATA[6]),
                      .MU1_EFPGA_MATHB_OPER_DATA_5_(MU1_EFPGA_MATHB_OPER_DATA[5]),
                      .MU1_EFPGA_MATHB_COEF_DATA_29_(MU1_EFPGA_MATHB_COEF_DATA[29]),
                      .MU1_EFPGA_MATHB_COEF_DATA_28_(MU1_EFPGA_MATHB_COEF_DATA[28]),
                      .MU1_EFPGA_MATHB_COEF_DATA_27_(MU1_EFPGA_MATHB_COEF_DATA[27]),
                      .MU1_EFPGA_MATHB_COEF_DATA_26_(MU1_EFPGA_MATHB_COEF_DATA[26]),
                      .MU1_EFPGA_MATHB_COEF_DATA_25_(MU1_EFPGA_MATHB_COEF_DATA[25]),
                      .MU1_EFPGA_MATHB_COEF_DATA_24_(MU1_EFPGA_MATHB_COEF_DATA[24]),
                      .MU1_EFPGA_MATHB_COEF_DATA_23_(MU1_EFPGA_MATHB_COEF_DATA[23]),
                      .MU1_EFPGA_MATHB_COEF_DATA_22_(MU1_EFPGA_MATHB_COEF_DATA[22]),
                      .MU1_EFPGA_MATHB_OPER_DATA_4_(MU1_EFPGA_MATHB_OPER_DATA[4]),
                      .MU1_EFPGA_MATHB_OPER_DATA_3_(MU1_EFPGA_MATHB_OPER_DATA[3]),
                      .MU1_EFPGA_MATHB_OPER_DATA_2_(MU1_EFPGA_MATHB_OPER_DATA[2]),
                      .MU1_EFPGA_MATHB_OPER_DATA_1_(MU1_EFPGA_MATHB_OPER_DATA[1]),
                      .MU1_EFPGA_MATHB_OPER_DATA_0_(MU1_EFPGA_MATHB_OPER_DATA[0]),
                      .MU1_EFPGA_MATHB_COEF_SEL(MU1_EFPGA_MATHB_COEF_SEL),
                      .MU1_EFPGA_MATHB_COEF_DATA_31_(MU1_EFPGA_MATHB_COEF_DATA[31]),
                      .MU1_EFPGA_MATHB_COEF_DATA_30_(MU1_EFPGA_MATHB_COEF_DATA[30]),
                      .MU1_EFPGA_MATHB_COEF_DATA_21_(MU1_EFPGA_MATHB_COEF_DATA[21]),
                      .MU1_EFPGA_MATHB_COEF_DATA_20_(MU1_EFPGA_MATHB_COEF_DATA[20]),
                      .MU1_EFPGA_MATHB_COEF_DATA_11_(MU1_EFPGA_MATHB_COEF_DATA[11]),
                      .MU1_EFPGA_MATHB_COEF_DATA_10_(MU1_EFPGA_MATHB_COEF_DATA[10]),
                      .MU1_EFPGA_MATHB_COEF_DATA_19_(MU1_EFPGA_MATHB_COEF_DATA[19]),
                      .MU1_EFPGA_MATHB_COEF_DATA_18_(MU1_EFPGA_MATHB_COEF_DATA[18]),
                      .MU1_EFPGA_MATHB_COEF_DATA_17_(MU1_EFPGA_MATHB_COEF_DATA[17]),
                      .MU1_EFPGA_MATHB_COEF_DATA_16_(MU1_EFPGA_MATHB_COEF_DATA[16]),
                      .MU1_EFPGA_MATHB_COEF_DATA_15_(MU1_EFPGA_MATHB_COEF_DATA[15]),
                      .MU1_EFPGA_MATHB_COEF_DATA_14_(MU1_EFPGA_MATHB_COEF_DATA[14]),
                      .MU1_EFPGA_MATHB_COEF_DATA_13_(MU1_EFPGA_MATHB_COEF_DATA[13]),
                      .MU1_EFPGA_MATHB_COEF_DATA_12_(MU1_EFPGA_MATHB_COEF_DATA[12]),
                      .MU1_EFPGA_MATHB_COEF_DATA_9_(MU1_EFPGA_MATHB_COEF_DATA[9]),
                      .MU1_EFPGA_MATHB_COEF_DATA_8_(MU1_EFPGA_MATHB_COEF_DATA[8]),
                      .MU1_EFPGA_MATHB_DATAOUT_SEL_1_(MU1_EFPGA_MATHB_DATAOUT_SEL[1]),
                      .MU1_EFPGA_MATHB_DATAOUT_SEL_0_(MU1_EFPGA_MATHB_DATAOUT_SEL[0]),
                      .MU1_EFPGA_TPRAM_COEF_W_MODE_1_(MU1_EFPGA_TPRAM_COEF_W_MODE[1]),
                      .MU1_EFPGA_TPRAM_COEF_W_MODE_0_(MU1_EFPGA_TPRAM_COEF_W_MODE[0]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_31_(MU1_EFPGA_TPRAM_COEF_W_DATA[31]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_30_(MU1_EFPGA_TPRAM_COEF_W_DATA[30]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_29_(MU1_EFPGA_TPRAM_COEF_W_DATA[29]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_28_(MU1_EFPGA_TPRAM_COEF_W_DATA[28]),
                      .MU1_EFPGA_MATHB_COEF_DATA_7_(MU1_EFPGA_MATHB_COEF_DATA[7]),
                      .MU1_EFPGA_MATHB_COEF_DATA_6_(MU1_EFPGA_MATHB_COEF_DATA[6]),
                      .MU1_EFPGA_MATHB_COEF_DATA_5_(MU1_EFPGA_MATHB_COEF_DATA[5]),
                      .MU1_EFPGA_MATHB_COEF_DATA_4_(MU1_EFPGA_MATHB_COEF_DATA[4]),
                      .MU1_EFPGA_MATHB_COEF_DATA_3_(MU1_EFPGA_MATHB_COEF_DATA[3]),
                      .MU1_EFPGA_MATHB_COEF_DATA_2_(MU1_EFPGA_MATHB_COEF_DATA[2]),
                      .MU1_EFPGA_MATHB_COEF_DATA_1_(MU1_EFPGA_MATHB_COEF_DATA[1]),
                      .MU1_EFPGA_MATHB_COEF_DATA_0_(MU1_EFPGA_MATHB_COEF_DATA[0]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_27_(MU1_EFPGA_TPRAM_COEF_W_DATA[27]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_26_(MU1_EFPGA_TPRAM_COEF_W_DATA[26]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_17_(MU1_EFPGA_TPRAM_COEF_W_DATA[17]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_16_(MU1_EFPGA_TPRAM_COEF_W_DATA[16]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_25_(MU1_EFPGA_TPRAM_COEF_W_DATA[25]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_24_(MU1_EFPGA_TPRAM_COEF_W_DATA[24]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_23_(MU1_EFPGA_TPRAM_COEF_W_DATA[23]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_22_(MU1_EFPGA_TPRAM_COEF_W_DATA[22]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_21_(MU1_EFPGA_TPRAM_COEF_W_DATA[21]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_20_(MU1_EFPGA_TPRAM_COEF_W_DATA[20]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_19_(MU1_EFPGA_TPRAM_COEF_W_DATA[19]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_18_(MU1_EFPGA_TPRAM_COEF_W_DATA[18]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_15_(MU1_EFPGA_TPRAM_COEF_W_DATA[15]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_14_(MU1_EFPGA_TPRAM_COEF_W_DATA[14]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_5_(MU1_EFPGA_TPRAM_COEF_W_DATA[5]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_4_(MU1_EFPGA_TPRAM_COEF_W_DATA[4]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_3_(MU1_EFPGA_TPRAM_COEF_W_DATA[3]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_2_(MU1_EFPGA_TPRAM_COEF_W_DATA[2]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_1_(MU1_EFPGA_TPRAM_COEF_W_DATA[1]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_0_(MU1_EFPGA_TPRAM_COEF_W_DATA[0]),
                      .MU1_EFPGA_TPRAM_COEF_W_CLK(MU1_EFPGA_TPRAM_COEF_W_CLK),
                      .MU1_EFPGA_TPRAM_COEF_W_ADDR_11_(MU1_EFPGA_TPRAM_COEF_W_ADDR[11]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_13_(MU1_EFPGA_TPRAM_COEF_W_DATA[13]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_12_(MU1_EFPGA_TPRAM_COEF_W_DATA[12]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_11_(MU1_EFPGA_TPRAM_COEF_W_DATA[11]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_10_(MU1_EFPGA_TPRAM_COEF_W_DATA[10]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_9_(MU1_EFPGA_TPRAM_COEF_W_DATA[9]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_8_(MU1_EFPGA_TPRAM_COEF_W_DATA[8]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_7_(MU1_EFPGA_TPRAM_COEF_W_DATA[7]),
                      .MU1_EFPGA_TPRAM_COEF_W_DATA_6_(MU1_EFPGA_TPRAM_COEF_W_DATA[6]),
                      .MU1_EFPGA_TPRAM_COEF_W_ADDR_10_(MU1_EFPGA_TPRAM_COEF_W_ADDR[10]),
                      .MU1_EFPGA_TPRAM_COEF_W_ADDR_9_(MU1_EFPGA_TPRAM_COEF_W_ADDR[9]),
                      .MU1_EFPGA_TPRAM_COEF_W_ADDR_0_(MU1_EFPGA_TPRAM_COEF_W_ADDR[0]),
                      .MU1_EFPGA_TPRAM_COEF_WE(MU1_EFPGA_TPRAM_COEF_WE),
                      .MU1_EFPGA_TPRAM_COEF_W_ADDR_8_(MU1_EFPGA_TPRAM_COEF_W_ADDR[8]),
                      .MU1_EFPGA_TPRAM_COEF_W_ADDR_7_(MU1_EFPGA_TPRAM_COEF_W_ADDR[7]),
                      .MU1_EFPGA_TPRAM_COEF_W_ADDR_6_(MU1_EFPGA_TPRAM_COEF_W_ADDR[6]),
                      .MU1_EFPGA_TPRAM_COEF_W_ADDR_5_(MU1_EFPGA_TPRAM_COEF_W_ADDR[5]),
                      .MU1_EFPGA_TPRAM_COEF_W_ADDR_4_(MU1_EFPGA_TPRAM_COEF_W_ADDR[4]),
                      .MU1_EFPGA_TPRAM_COEF_W_ADDR_3_(MU1_EFPGA_TPRAM_COEF_W_ADDR[3]),
                      .MU1_EFPGA_TPRAM_COEF_W_ADDR_2_(MU1_EFPGA_TPRAM_COEF_W_ADDR[2]),
                      .MU1_EFPGA_TPRAM_COEF_W_ADDR_1_(MU1_EFPGA_TPRAM_COEF_W_ADDR[1]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_25_(MU0_EFPGA_TPRAM_OPER_W_DATA[25]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_24_(MU0_EFPGA_TPRAM_OPER_W_DATA[24]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_23_(MU0_EFPGA_TPRAM_OPER_W_DATA[23]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_22_(MU0_EFPGA_TPRAM_OPER_W_DATA[22]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_21_(MU0_EFPGA_TPRAM_OPER_W_DATA[21]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_20_(MU0_EFPGA_TPRAM_OPER_W_DATA[20]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_19_(MU0_EFPGA_TPRAM_OPER_W_DATA[19]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_18_(MU0_EFPGA_TPRAM_OPER_W_DATA[18]),
                      .MU0_EFPGA_TPRAM_OPER_W_MODE_1_(MU0_EFPGA_TPRAM_OPER_W_MODE[1]),
                      .MU0_EFPGA_TPRAM_OPER_W_MODE_0_(MU0_EFPGA_TPRAM_OPER_W_MODE[0]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_31_(MU0_EFPGA_TPRAM_OPER_W_DATA[31]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_30_(MU0_EFPGA_TPRAM_OPER_W_DATA[30]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_29_(MU0_EFPGA_TPRAM_OPER_W_DATA[29]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_28_(MU0_EFPGA_TPRAM_OPER_W_DATA[28]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_27_(MU0_EFPGA_TPRAM_OPER_W_DATA[27]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_26_(MU0_EFPGA_TPRAM_OPER_W_DATA[26]),
                      .MU1_EFPGA_TPRAM_COEF_WDSEL(MU1_EFPGA_TPRAM_COEF_WDSEL),
                      .MU1_EFPGA_TPRAM_COEF_R_MODE_1_(MU1_EFPGA_TPRAM_COEF_R_MODE[1]),
                      .MU1_EFPGA_TPRAM_COEF_R_ADDR_5_(MU1_EFPGA_TPRAM_COEF_R_ADDR[5]),
                      .MU1_EFPGA_TPRAM_COEF_R_ADDR_4_(MU1_EFPGA_TPRAM_COEF_R_ADDR[4]),
                      .MU1_EFPGA_TPRAM_COEF_R_ADDR_3_(MU1_EFPGA_TPRAM_COEF_R_ADDR[3]),
                      .MU1_EFPGA_TPRAM_COEF_R_ADDR_2_(MU1_EFPGA_TPRAM_COEF_R_ADDR[2]),
                      .MU1_EFPGA_TPRAM_COEF_R_ADDR_1_(MU1_EFPGA_TPRAM_COEF_R_ADDR[1]),
                      .MU1_EFPGA_TPRAM_COEF_R_ADDR_0_(MU1_EFPGA_TPRAM_COEF_R_ADDR[0]),
                      .MU1_EFPGA_TPRAM_COEF_POWERDN(MU1_EFPGA_TPRAM_COEF_POWERDN),
                      .MU1_EFPGA_TPRAM_COEF_R_MODE_0_(MU1_EFPGA_TPRAM_COEF_R_MODE[0]),
                      .MU1_EFPGA_TPRAM_COEF_R_CLK(MU1_EFPGA_TPRAM_COEF_R_CLK),
                      .MU1_EFPGA_TPRAM_COEF_R_ADDR_11_(MU1_EFPGA_TPRAM_COEF_R_ADDR[11]),
                      .MU1_EFPGA_TPRAM_COEF_R_ADDR_10_(MU1_EFPGA_TPRAM_COEF_R_ADDR[10]),
                      .MU1_EFPGA_TPRAM_COEF_R_ADDR_9_(MU1_EFPGA_TPRAM_COEF_R_ADDR[9]),
                      .MU1_EFPGA_TPRAM_COEF_R_ADDR_8_(MU1_EFPGA_TPRAM_COEF_R_ADDR[8]),
                      .MU1_EFPGA_TPRAM_COEF_R_ADDR_7_(MU1_EFPGA_TPRAM_COEF_R_ADDR[7]),
                      .MU1_EFPGA_TPRAM_COEF_R_ADDR_6_(MU1_EFPGA_TPRAM_COEF_R_ADDR[6]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_17_(MU0_EFPGA_TPRAM_OPER_W_DATA[17]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_16_(MU0_EFPGA_TPRAM_OPER_W_DATA[16]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_7_(MU0_EFPGA_TPRAM_OPER_W_DATA[7]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_6_(MU0_EFPGA_TPRAM_OPER_W_DATA[6]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_15_(MU0_EFPGA_TPRAM_OPER_W_DATA[15]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_14_(MU0_EFPGA_TPRAM_OPER_W_DATA[14]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_13_(MU0_EFPGA_TPRAM_OPER_W_DATA[13]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_12_(MU0_EFPGA_TPRAM_OPER_W_DATA[12]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_11_(MU0_EFPGA_TPRAM_OPER_W_DATA[11]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_10_(MU0_EFPGA_TPRAM_OPER_W_DATA[10]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_9_(MU0_EFPGA_TPRAM_OPER_W_DATA[9]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_8_(MU0_EFPGA_TPRAM_OPER_W_DATA[8]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_5_(MU0_EFPGA_TPRAM_OPER_W_DATA[5]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_4_(MU0_EFPGA_TPRAM_OPER_W_DATA[4]),
                      .MU0_EFPGA_TPRAM_OPER_W_ADDR_8_(MU0_EFPGA_TPRAM_OPER_W_ADDR[8]),
                      .MU0_EFPGA_TPRAM_OPER_W_ADDR_7_(MU0_EFPGA_TPRAM_OPER_W_ADDR[7]),
                      .MU0_EFPGA_TPRAM_OPER_W_ADDR_6_(MU0_EFPGA_TPRAM_OPER_W_ADDR[6]),
                      .MU0_EFPGA_TPRAM_OPER_W_ADDR_5_(MU0_EFPGA_TPRAM_OPER_W_ADDR[5]),
                      .MU0_EFPGA_TPRAM_OPER_W_ADDR_4_(MU0_EFPGA_TPRAM_OPER_W_ADDR[4]),
                      .MU0_EFPGA_TPRAM_OPER_W_ADDR_3_(MU0_EFPGA_TPRAM_OPER_W_ADDR[3]),
                      .MU0_EFPGA_TPRAM_OPER_W_ADDR_2_(MU0_EFPGA_TPRAM_OPER_W_ADDR[2]),
                      .MU0_EFPGA_TPRAM_OPER_W_ADDR_1_(MU0_EFPGA_TPRAM_OPER_W_ADDR[1]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_3_(MU0_EFPGA_TPRAM_OPER_W_DATA[3]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_2_(MU0_EFPGA_TPRAM_OPER_W_DATA[2]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_1_(MU0_EFPGA_TPRAM_OPER_W_DATA[1]),
                      .MU0_EFPGA_TPRAM_OPER_W_DATA_0_(MU0_EFPGA_TPRAM_OPER_W_DATA[0]),
                      .MU0_EFPGA_TPRAM_OPER_W_CLK(MU0_EFPGA_TPRAM_OPER_W_CLK),
                      .MU0_EFPGA_TPRAM_OPER_W_ADDR_11_(MU0_EFPGA_TPRAM_OPER_W_ADDR[11]),
                      .MU0_EFPGA_TPRAM_OPER_W_ADDR_10_(MU0_EFPGA_TPRAM_OPER_W_ADDR[10]),
                      .MU0_EFPGA_TPRAM_OPER_W_ADDR_9_(MU0_EFPGA_TPRAM_OPER_W_ADDR[9]),
                      .MU0_EFPGA_TPRAM_OPER_W_ADDR_0_(MU0_EFPGA_TPRAM_OPER_W_ADDR[0]),
                      .MU0_EFPGA_TPRAM_OPER_WE(MU0_EFPGA_TPRAM_OPER_WE),
                      .MU0_EFPGA_TPRAM_OPER_R_ADDR_7_(MU0_EFPGA_TPRAM_OPER_R_ADDR[7]),
                      .MU0_EFPGA_TPRAM_OPER_R_ADDR_6_(MU0_EFPGA_TPRAM_OPER_R_ADDR[6]),
                      .MU0_EFPGA_TPRAM_OPER_WDSEL(MU0_EFPGA_TPRAM_OPER_WDSEL),
                      .MU0_EFPGA_TPRAM_OPER_R_MODE_1_(MU0_EFPGA_TPRAM_OPER_R_MODE[1]),
                      .MU0_EFPGA_TPRAM_OPER_R_MODE_0_(MU0_EFPGA_TPRAM_OPER_R_MODE[0]),
                      .MU0_EFPGA_TPRAM_OPER_R_CLK(MU0_EFPGA_TPRAM_OPER_R_CLK),
                      .MU0_EFPGA_TPRAM_OPER_R_ADDR_11_(MU0_EFPGA_TPRAM_OPER_R_ADDR[11]),
                      .MU0_EFPGA_TPRAM_OPER_R_ADDR_10_(MU0_EFPGA_TPRAM_OPER_R_ADDR[10]),
                      .MU0_EFPGA_TPRAM_OPER_R_ADDR_9_(MU0_EFPGA_TPRAM_OPER_R_ADDR[9]),
                      .MU0_EFPGA_TPRAM_OPER_R_ADDR_8_(MU0_EFPGA_TPRAM_OPER_R_ADDR[8]),
                      .MU0_EFPGA_TPRAM_OPER_R_ADDR_5_(MU0_EFPGA_TPRAM_OPER_R_ADDR[5]),
                      .MU0_EFPGA_TPRAM_OPER_R_ADDR_4_(MU0_EFPGA_TPRAM_OPER_R_ADDR[4]),
                      .MU0_EFPGA_MATHB_MAC_OUT_SEL_4_(MU0_EFPGA_MATHB_MAC_OUT_SEL[4]),
                      .MU0_EFPGA_MATHB_MAC_OUT_SEL_3_(MU0_EFPGA_MATHB_MAC_OUT_SEL[3]),
                      .MU0_EFPGA_MATHB_MAC_OUT_SEL_2_(MU0_EFPGA_MATHB_MAC_OUT_SEL[2]),
                      .MU0_EFPGA_MATHB_MAC_OUT_SEL_1_(MU0_EFPGA_MATHB_MAC_OUT_SEL[1]),
                      .MU0_EFPGA_MATHB_MAC_OUT_SEL_0_(MU0_EFPGA_MATHB_MAC_OUT_SEL[0]),
                      .MU0_EFPGA_MATHB_MAC_ACC_SAT(MU0_EFPGA_MATHB_MAC_ACC_SAT),
                      .MU0_EFPGA_MATHB_MAC_ACC_RND(MU0_EFPGA_MATHB_MAC_ACC_RND),
                      .MU0_EFPGA_MATHB_MAC_ACC_CLEAR(MU0_EFPGA_MATHB_MAC_ACC_CLEAR),
                      .MU0_EFPGA_TPRAM_OPER_R_ADDR_3_(MU0_EFPGA_TPRAM_OPER_R_ADDR[3]),
                      .MU0_EFPGA_TPRAM_OPER_R_ADDR_2_(MU0_EFPGA_TPRAM_OPER_R_ADDR[2]),
                      .MU0_EFPGA_TPRAM_OPER_R_ADDR_1_(MU0_EFPGA_TPRAM_OPER_R_ADDR[1]),
                      .MU0_EFPGA_TPRAM_OPER_R_ADDR_0_(MU0_EFPGA_TPRAM_OPER_R_ADDR[0]),
                      .MU0_EFPGA_TPRAM_OPER_POWERDN(MU0_EFPGA_TPRAM_OPER_POWERDN),
                      .MU0_EFPGA2MATHB_CLK(MU0_EFPGA2MATHB_CLK),
                      .MU0_EFPGA_MATHB_CLK_EN(MU0_EFPGA_MATHB_CLK_EN),
                      .MU0_EFPGA_MATHB_MAC_OUT_SEL_5_(MU0_EFPGA_MATHB_MAC_OUT_SEL[5]),
                      .MU0_EFPGA_MATHB_OPER_SEL(MU0_EFPGA_MATHB_OPER_SEL),
                      .MU0_EFPGA_MATHB_OPER_DATA_31_(MU0_EFPGA_MATHB_OPER_DATA[31]),
                      .MU0_EFPGA_MATHB_OPER_DATA_22_(MU0_EFPGA_MATHB_OPER_DATA[22]),
                      .MU0_EFPGA_MATHB_OPER_DATA_21_(MU0_EFPGA_MATHB_OPER_DATA[21]),
                      .MU0_EFPGA_MATHB_OPER_DATA_30_(MU0_EFPGA_MATHB_OPER_DATA[30]),
                      .MU0_EFPGA_MATHB_OPER_DATA_29_(MU0_EFPGA_MATHB_OPER_DATA[29]),
                      .MU0_EFPGA_MATHB_OPER_DATA_28_(MU0_EFPGA_MATHB_OPER_DATA[28]),
                      .MU0_EFPGA_MATHB_OPER_DATA_27_(MU0_EFPGA_MATHB_OPER_DATA[27]),
                      .MU0_EFPGA_MATHB_OPER_DATA_26_(MU0_EFPGA_MATHB_OPER_DATA[26]),
                      .MU0_EFPGA_MATHB_OPER_DATA_25_(MU0_EFPGA_MATHB_OPER_DATA[25]),
                      .MU0_EFPGA_MATHB_OPER_DATA_24_(MU0_EFPGA_MATHB_OPER_DATA[24]),
                      .MU0_EFPGA_MATHB_OPER_DATA_23_(MU0_EFPGA_MATHB_OPER_DATA[23]),
                      .MU0_EFPGA_MATHB_OPER_DATA_20_(MU0_EFPGA_MATHB_OPER_DATA[20]),
                      .MU0_EFPGA_MATHB_OPER_DATA_19_(MU0_EFPGA_MATHB_OPER_DATA[19]),
                      .MU0_EFPGA_MATHB_OPER_DATA_10_(MU0_EFPGA_MATHB_OPER_DATA[10]),
                      .MU0_EFPGA_MATHB_OPER_DATA_9_(MU0_EFPGA_MATHB_OPER_DATA[9]),
                      .MU0_EFPGA_MATHB_OPER_DATA_8_(MU0_EFPGA_MATHB_OPER_DATA[8]),
                      .MU0_EFPGA_MATHB_OPER_DATA_7_(MU0_EFPGA_MATHB_OPER_DATA[7]),
                      .MU0_EFPGA_MATHB_OPER_DATA_6_(MU0_EFPGA_MATHB_OPER_DATA[6]),
                      .MU0_EFPGA_MATHB_OPER_DATA_5_(MU0_EFPGA_MATHB_OPER_DATA[5]),
                      .MU0_EFPGA_MATHB_OPER_DATA_4_(MU0_EFPGA_MATHB_OPER_DATA[4]),
                      .MU0_EFPGA_MATHB_OPER_DATA_3_(MU0_EFPGA_MATHB_OPER_DATA[3]),
                      .MU0_EFPGA_MATHB_OPER_DATA_18_(MU0_EFPGA_MATHB_OPER_DATA[18]),
                      .MU0_EFPGA_MATHB_OPER_DATA_17_(MU0_EFPGA_MATHB_OPER_DATA[17]),
                      .MU0_EFPGA_MATHB_OPER_DATA_16_(MU0_EFPGA_MATHB_OPER_DATA[16]),
                      .MU0_EFPGA_MATHB_OPER_DATA_15_(MU0_EFPGA_MATHB_OPER_DATA[15]),
                      .MU0_EFPGA_MATHB_OPER_DATA_14_(MU0_EFPGA_MATHB_OPER_DATA[14]),
                      .MU0_EFPGA_MATHB_OPER_DATA_13_(MU0_EFPGA_MATHB_OPER_DATA[13]),
                      .MU0_EFPGA_MATHB_OPER_DATA_12_(MU0_EFPGA_MATHB_OPER_DATA[12]),
                      .MU0_EFPGA_MATHB_OPER_DATA_11_(MU0_EFPGA_MATHB_OPER_DATA[11]),
                      .MU0_EFPGA_MATHB_OPER_DATA_2_(MU0_EFPGA_MATHB_OPER_DATA[2]),
                      .MU0_EFPGA_MATHB_OPER_DATA_1_(MU0_EFPGA_MATHB_OPER_DATA[1]),
                      .MU0_EFPGA_MATHB_COEF_DATA_25_(MU0_EFPGA_MATHB_COEF_DATA[25]),
                      .MU0_EFPGA_MATHB_COEF_DATA_24_(MU0_EFPGA_MATHB_COEF_DATA[24]),
                      .MU0_EFPGA_MATHB_OPER_DATA_0_(MU0_EFPGA_MATHB_OPER_DATA[0]),
                      .MU0_EFPGA_MATHB_COEF_SEL(MU0_EFPGA_MATHB_COEF_SEL),
                      .MU0_EFPGA_MATHB_COEF_DATA_31_(MU0_EFPGA_MATHB_COEF_DATA[31]),
                      .MU0_EFPGA_MATHB_COEF_DATA_30_(MU0_EFPGA_MATHB_COEF_DATA[30]),
                      .MU0_EFPGA_MATHB_COEF_DATA_29_(MU0_EFPGA_MATHB_COEF_DATA[29]),
                      .MU0_EFPGA_MATHB_COEF_DATA_28_(MU0_EFPGA_MATHB_COEF_DATA[28]),
                      .MU0_EFPGA_MATHB_COEF_DATA_27_(MU0_EFPGA_MATHB_COEF_DATA[27]),
                      .MU0_EFPGA_MATHB_COEF_DATA_26_(MU0_EFPGA_MATHB_COEF_DATA[26]),
                      .MU1_EFPGA_MATHB_TC_defPin(MU1_EFPGA_MATHB_TC_defPin),
                      .MU1_EFPGA_MATHB_OPER_defPin_1_(MU1_EFPGA_MATHB_OPER_defPin[1]),
                      .MU1_EFPGA_MATHB_OPER_defPin_0_(MU1_EFPGA_MATHB_OPER_defPin[0]),
                      .MU1_EFPGA_MATHB_COEF_defPin_1_(MU1_EFPGA_MATHB_COEF_defPin[1]),
                      .MU1_EFPGA_MATHB_COEF_defPin_0_(MU1_EFPGA_MATHB_COEF_defPin[0]),
                      .MU0_EFPGA_MATHB_TC_defPin(MU0_EFPGA_MATHB_TC_defPin),
                      .MU0_EFPGA_MATHB_OPER_defPin_1_(MU0_EFPGA_MATHB_OPER_defPin[1]),
                      .MU0_EFPGA_MATHB_OPER_defPin_0_(MU0_EFPGA_MATHB_OPER_defPin[0]),
                      .MU0_EFPGA_MATHB_COEF_defPin_1_(MU0_EFPGA_MATHB_COEF_defPin[1]),
                      .MU0_EFPGA_MATHB_COEF_defPin_0_(MU0_EFPGA_MATHB_COEF_defPin[0]),

                      // Inputs
                      .MU0_MATHB_EFPGA_MAC_OUT_7_(MU0_MATHB_EFPGA_MAC_OUT[7]),
                      .MU0_MATHB_EFPGA_MAC_OUT_6_(MU0_MATHB_EFPGA_MAC_OUT[6]),
                      .MU0_MATHB_EFPGA_MAC_OUT_5_(MU0_MATHB_EFPGA_MAC_OUT[5]),
                      .MU0_MATHB_EFPGA_MAC_OUT_4_(MU0_MATHB_EFPGA_MAC_OUT[4]),
                      .MU0_MATHB_EFPGA_MAC_OUT_3_(MU0_MATHB_EFPGA_MAC_OUT[3]),
                      .MU0_MATHB_EFPGA_MAC_OUT_2_(MU0_MATHB_EFPGA_MAC_OUT[2]),
                      .MU0_MATHB_EFPGA_MAC_OUT_1_(MU0_MATHB_EFPGA_MAC_OUT[1]),
                      .MU0_MATHB_EFPGA_MAC_OUT_0_(MU0_MATHB_EFPGA_MAC_OUT[0]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_31_(MU0_TPRAM_EFPGA_COEF_R_DATA[31]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_30_(MU0_TPRAM_EFPGA_COEF_R_DATA[30]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_29_(MU0_TPRAM_EFPGA_COEF_R_DATA[29]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_28_(MU0_TPRAM_EFPGA_COEF_R_DATA[28]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_27_(MU0_TPRAM_EFPGA_COEF_R_DATA[27]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_26_(MU0_TPRAM_EFPGA_COEF_R_DATA[26]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_25_(MU0_TPRAM_EFPGA_COEF_R_DATA[25]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_24_(MU0_TPRAM_EFPGA_COEF_R_DATA[24]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_23_(MU0_TPRAM_EFPGA_COEF_R_DATA[23]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_22_(MU0_TPRAM_EFPGA_COEF_R_DATA[22]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_21_(MU0_TPRAM_EFPGA_COEF_R_DATA[21]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_20_(MU0_TPRAM_EFPGA_COEF_R_DATA[20]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_19_(MU0_TPRAM_EFPGA_COEF_R_DATA[19]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_18_(MU0_TPRAM_EFPGA_COEF_R_DATA[18]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_17_(MU0_TPRAM_EFPGA_COEF_R_DATA[17]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_16_(MU0_TPRAM_EFPGA_COEF_R_DATA[16]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_15_(MU0_TPRAM_EFPGA_COEF_R_DATA[15]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_14_(MU0_TPRAM_EFPGA_COEF_R_DATA[14]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_13_(MU0_TPRAM_EFPGA_COEF_R_DATA[13]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_12_(MU0_TPRAM_EFPGA_COEF_R_DATA[12]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_11_(MU0_TPRAM_EFPGA_COEF_R_DATA[11]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_10_(MU0_TPRAM_EFPGA_COEF_R_DATA[10]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_9_(MU0_TPRAM_EFPGA_COEF_R_DATA[9]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_8_(MU0_TPRAM_EFPGA_COEF_R_DATA[8]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_7_(MU0_TPRAM_EFPGA_COEF_R_DATA[7]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_6_(MU0_TPRAM_EFPGA_COEF_R_DATA[6]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_5_(MU0_TPRAM_EFPGA_COEF_R_DATA[5]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_4_(MU0_TPRAM_EFPGA_COEF_R_DATA[4]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_3_(MU0_TPRAM_EFPGA_COEF_R_DATA[3]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_2_(MU0_TPRAM_EFPGA_COEF_R_DATA[2]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_1_(MU0_TPRAM_EFPGA_COEF_R_DATA[1]),
                      .MU0_TPRAM_EFPGA_COEF_R_DATA_0_(MU0_TPRAM_EFPGA_COEF_R_DATA[0]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_31_(MU1_TPRAM_EFPGA_OPER_R_DATA[31]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_30_(MU1_TPRAM_EFPGA_OPER_R_DATA[30]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_29_(MU1_TPRAM_EFPGA_OPER_R_DATA[29]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_28_(MU1_TPRAM_EFPGA_OPER_R_DATA[28]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_27_(MU1_TPRAM_EFPGA_OPER_R_DATA[27]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_26_(MU1_TPRAM_EFPGA_OPER_R_DATA[26]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_25_(MU1_TPRAM_EFPGA_OPER_R_DATA[25]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_24_(MU1_TPRAM_EFPGA_OPER_R_DATA[24]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_23_(MU1_TPRAM_EFPGA_OPER_R_DATA[23]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_22_(MU1_TPRAM_EFPGA_OPER_R_DATA[22]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_21_(MU1_TPRAM_EFPGA_OPER_R_DATA[21]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_20_(MU1_TPRAM_EFPGA_OPER_R_DATA[20]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_19_(MU1_TPRAM_EFPGA_OPER_R_DATA[19]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_18_(MU1_TPRAM_EFPGA_OPER_R_DATA[18]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_17_(MU1_TPRAM_EFPGA_OPER_R_DATA[17]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_16_(MU1_TPRAM_EFPGA_OPER_R_DATA[16]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_15_(MU1_TPRAM_EFPGA_OPER_R_DATA[15]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_14_(MU1_TPRAM_EFPGA_OPER_R_DATA[14]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_13_(MU1_TPRAM_EFPGA_OPER_R_DATA[13]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_12_(MU1_TPRAM_EFPGA_OPER_R_DATA[12]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_31_(MU0_TPRAM_EFPGA_OPER_R_DATA[31]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_30_(MU0_TPRAM_EFPGA_OPER_R_DATA[30]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_29_(MU0_TPRAM_EFPGA_OPER_R_DATA[29]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_28_(MU0_TPRAM_EFPGA_OPER_R_DATA[28]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_11_(MU1_TPRAM_EFPGA_OPER_R_DATA[11]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_10_(MU1_TPRAM_EFPGA_OPER_R_DATA[10]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_9_(MU1_TPRAM_EFPGA_OPER_R_DATA[9]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_8_(MU1_TPRAM_EFPGA_OPER_R_DATA[8]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_7_(MU1_TPRAM_EFPGA_OPER_R_DATA[7]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_6_(MU1_TPRAM_EFPGA_OPER_R_DATA[6]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_5_(MU1_TPRAM_EFPGA_OPER_R_DATA[5]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_4_(MU1_TPRAM_EFPGA_OPER_R_DATA[4]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_3_(MU1_TPRAM_EFPGA_OPER_R_DATA[3]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_2_(MU1_TPRAM_EFPGA_OPER_R_DATA[2]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_1_(MU1_TPRAM_EFPGA_OPER_R_DATA[1]),
                      .MU1_TPRAM_EFPGA_OPER_R_DATA_0_(MU1_TPRAM_EFPGA_OPER_R_DATA[0]),
                      .MU1_MATHB_EFPGA_MAC_OUT_31_(MU1_MATHB_EFPGA_MAC_OUT[31]),
                      .MU1_MATHB_EFPGA_MAC_OUT_30_(MU1_MATHB_EFPGA_MAC_OUT[30]),
                      .MU1_MATHB_EFPGA_MAC_OUT_29_(MU1_MATHB_EFPGA_MAC_OUT[29]),
                      .MU1_MATHB_EFPGA_MAC_OUT_28_(MU1_MATHB_EFPGA_MAC_OUT[28]),
                      .MU1_MATHB_EFPGA_MAC_OUT_27_(MU1_MATHB_EFPGA_MAC_OUT[27]),
                      .MU1_MATHB_EFPGA_MAC_OUT_26_(MU1_MATHB_EFPGA_MAC_OUT[26]),
                      .MU1_MATHB_EFPGA_MAC_OUT_25_(MU1_MATHB_EFPGA_MAC_OUT[25]),
                      .MU1_MATHB_EFPGA_MAC_OUT_24_(MU1_MATHB_EFPGA_MAC_OUT[24]),
                      .MU1_MATHB_EFPGA_MAC_OUT_23_(MU1_MATHB_EFPGA_MAC_OUT[23]),
                      .MU1_MATHB_EFPGA_MAC_OUT_22_(MU1_MATHB_EFPGA_MAC_OUT[22]),
                      .MU1_MATHB_EFPGA_MAC_OUT_21_(MU1_MATHB_EFPGA_MAC_OUT[21]),
                      .MU1_MATHB_EFPGA_MAC_OUT_20_(MU1_MATHB_EFPGA_MAC_OUT[20]),
                      .MU1_MATHB_EFPGA_MAC_OUT_19_(MU1_MATHB_EFPGA_MAC_OUT[19]),
                      .MU1_MATHB_EFPGA_MAC_OUT_18_(MU1_MATHB_EFPGA_MAC_OUT[18]),
                      .MU1_MATHB_EFPGA_MAC_OUT_17_(MU1_MATHB_EFPGA_MAC_OUT[17]),
                      .MU1_MATHB_EFPGA_MAC_OUT_16_(MU1_MATHB_EFPGA_MAC_OUT[16]),
                      .MU1_MATHB_EFPGA_MAC_OUT_15_(MU1_MATHB_EFPGA_MAC_OUT[15]),
                      .MU1_MATHB_EFPGA_MAC_OUT_14_(MU1_MATHB_EFPGA_MAC_OUT[14]),
                      .MU1_MATHB_EFPGA_MAC_OUT_13_(MU1_MATHB_EFPGA_MAC_OUT[13]),
                      .MU1_MATHB_EFPGA_MAC_OUT_12_(MU1_MATHB_EFPGA_MAC_OUT[12]),
                      .MU1_MATHB_EFPGA_MAC_OUT_11_(MU1_MATHB_EFPGA_MAC_OUT[11]),
                      .MU1_MATHB_EFPGA_MAC_OUT_10_(MU1_MATHB_EFPGA_MAC_OUT[10]),
                      .MU1_MATHB_EFPGA_MAC_OUT_9_(MU1_MATHB_EFPGA_MAC_OUT[9]),
                      .MU1_MATHB_EFPGA_MAC_OUT_8_(MU1_MATHB_EFPGA_MAC_OUT[8]),
                      .MU1_MATHB_EFPGA_MAC_OUT_7_(MU1_MATHB_EFPGA_MAC_OUT[7]),
                      .MU1_MATHB_EFPGA_MAC_OUT_6_(MU1_MATHB_EFPGA_MAC_OUT[6]),
                      .MU1_MATHB_EFPGA_MAC_OUT_5_(MU1_MATHB_EFPGA_MAC_OUT[5]),
                      .MU1_MATHB_EFPGA_MAC_OUT_4_(MU1_MATHB_EFPGA_MAC_OUT[4]),
                      .MU1_MATHB_EFPGA_MAC_OUT_3_(MU1_MATHB_EFPGA_MAC_OUT[3]),
                      .MU1_MATHB_EFPGA_MAC_OUT_2_(MU1_MATHB_EFPGA_MAC_OUT[2]),
                      .MU1_MATHB_EFPGA_MAC_OUT_1_(MU1_MATHB_EFPGA_MAC_OUT[1]),
                      .MU1_MATHB_EFPGA_MAC_OUT_0_(MU1_MATHB_EFPGA_MAC_OUT[0]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_31_(MU1_TPRAM_EFPGA_COEF_R_DATA[31]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_30_(MU1_TPRAM_EFPGA_COEF_R_DATA[30]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_29_(MU1_TPRAM_EFPGA_COEF_R_DATA[29]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_28_(MU1_TPRAM_EFPGA_COEF_R_DATA[28]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_27_(MU1_TPRAM_EFPGA_COEF_R_DATA[27]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_26_(MU1_TPRAM_EFPGA_COEF_R_DATA[26]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_25_(MU1_TPRAM_EFPGA_COEF_R_DATA[25]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_24_(MU1_TPRAM_EFPGA_COEF_R_DATA[24]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_23_(MU1_TPRAM_EFPGA_COEF_R_DATA[23]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_22_(MU1_TPRAM_EFPGA_COEF_R_DATA[22]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_21_(MU1_TPRAM_EFPGA_COEF_R_DATA[21]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_20_(MU1_TPRAM_EFPGA_COEF_R_DATA[20]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_19_(MU1_TPRAM_EFPGA_COEF_R_DATA[19]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_18_(MU1_TPRAM_EFPGA_COEF_R_DATA[18]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_27_(MU0_TPRAM_EFPGA_OPER_R_DATA[27]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_26_(MU0_TPRAM_EFPGA_OPER_R_DATA[26]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_25_(MU0_TPRAM_EFPGA_OPER_R_DATA[25]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_24_(MU0_TPRAM_EFPGA_OPER_R_DATA[24]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_23_(MU0_TPRAM_EFPGA_OPER_R_DATA[23]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_22_(MU0_TPRAM_EFPGA_OPER_R_DATA[22]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_21_(MU0_TPRAM_EFPGA_OPER_R_DATA[21]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_20_(MU0_TPRAM_EFPGA_OPER_R_DATA[20]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_17_(MU1_TPRAM_EFPGA_COEF_R_DATA[17]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_16_(MU1_TPRAM_EFPGA_COEF_R_DATA[16]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_15_(MU1_TPRAM_EFPGA_COEF_R_DATA[15]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_14_(MU1_TPRAM_EFPGA_COEF_R_DATA[14]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_13_(MU1_TPRAM_EFPGA_COEF_R_DATA[13]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_12_(MU1_TPRAM_EFPGA_COEF_R_DATA[12]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_11_(MU1_TPRAM_EFPGA_COEF_R_DATA[11]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_10_(MU1_TPRAM_EFPGA_COEF_R_DATA[10]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_9_(MU1_TPRAM_EFPGA_COEF_R_DATA[9]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_8_(MU1_TPRAM_EFPGA_COEF_R_DATA[8]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_7_(MU1_TPRAM_EFPGA_COEF_R_DATA[7]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_6_(MU1_TPRAM_EFPGA_COEF_R_DATA[6]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_5_(MU1_TPRAM_EFPGA_COEF_R_DATA[5]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_4_(MU1_TPRAM_EFPGA_COEF_R_DATA[4]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_3_(MU1_TPRAM_EFPGA_COEF_R_DATA[3]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_2_(MU1_TPRAM_EFPGA_COEF_R_DATA[2]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_1_(MU1_TPRAM_EFPGA_COEF_R_DATA[1]),
                      .MU1_TPRAM_EFPGA_COEF_R_DATA_0_(MU1_TPRAM_EFPGA_COEF_R_DATA[0]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_19_(MU0_TPRAM_EFPGA_OPER_R_DATA[19]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_18_(MU0_TPRAM_EFPGA_OPER_R_DATA[18]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_17_(MU0_TPRAM_EFPGA_OPER_R_DATA[17]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_16_(MU0_TPRAM_EFPGA_OPER_R_DATA[16]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_15_(MU0_TPRAM_EFPGA_OPER_R_DATA[15]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_14_(MU0_TPRAM_EFPGA_OPER_R_DATA[14]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_13_(MU0_TPRAM_EFPGA_OPER_R_DATA[13]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_12_(MU0_TPRAM_EFPGA_OPER_R_DATA[12]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_11_(MU0_TPRAM_EFPGA_OPER_R_DATA[11]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_10_(MU0_TPRAM_EFPGA_OPER_R_DATA[10]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_9_(MU0_TPRAM_EFPGA_OPER_R_DATA[9]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_8_(MU0_TPRAM_EFPGA_OPER_R_DATA[8]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_7_(MU0_TPRAM_EFPGA_OPER_R_DATA[7]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_6_(MU0_TPRAM_EFPGA_OPER_R_DATA[6]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_5_(MU0_TPRAM_EFPGA_OPER_R_DATA[5]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_4_(MU0_TPRAM_EFPGA_OPER_R_DATA[4]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_3_(MU0_TPRAM_EFPGA_OPER_R_DATA[3]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_2_(MU0_TPRAM_EFPGA_OPER_R_DATA[2]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_1_(MU0_TPRAM_EFPGA_OPER_R_DATA[1]),
                      .MU0_TPRAM_EFPGA_OPER_R_DATA_0_(MU0_TPRAM_EFPGA_OPER_R_DATA[0]),
                      .MU0_MATHB_EFPGA_MAC_OUT_31_(MU0_MATHB_EFPGA_MAC_OUT[31]),
                      .MU0_MATHB_EFPGA_MAC_OUT_30_(MU0_MATHB_EFPGA_MAC_OUT[30]),
                      .MU0_MATHB_EFPGA_MAC_OUT_29_(MU0_MATHB_EFPGA_MAC_OUT[29]),
                      .MU0_MATHB_EFPGA_MAC_OUT_28_(MU0_MATHB_EFPGA_MAC_OUT[28]),
                      .MU0_MATHB_EFPGA_MAC_OUT_27_(MU0_MATHB_EFPGA_MAC_OUT[27]),
                      .MU0_MATHB_EFPGA_MAC_OUT_26_(MU0_MATHB_EFPGA_MAC_OUT[26]),
                      .MU0_MATHB_EFPGA_MAC_OUT_25_(MU0_MATHB_EFPGA_MAC_OUT[25]),
                      .MU0_MATHB_EFPGA_MAC_OUT_24_(MU0_MATHB_EFPGA_MAC_OUT[24]),
                      .MU0_MATHB_EFPGA_MAC_OUT_23_(MU0_MATHB_EFPGA_MAC_OUT[23]),
                      .MU0_MATHB_EFPGA_MAC_OUT_22_(MU0_MATHB_EFPGA_MAC_OUT[22]),
                      .MU0_MATHB_EFPGA_MAC_OUT_21_(MU0_MATHB_EFPGA_MAC_OUT[21]),
                      .MU0_MATHB_EFPGA_MAC_OUT_20_(MU0_MATHB_EFPGA_MAC_OUT[20]),
                      .MU0_MATHB_EFPGA_MAC_OUT_19_(MU0_MATHB_EFPGA_MAC_OUT[19]),
                      .MU0_MATHB_EFPGA_MAC_OUT_18_(MU0_MATHB_EFPGA_MAC_OUT[18]),
                      .MU0_MATHB_EFPGA_MAC_OUT_17_(MU0_MATHB_EFPGA_MAC_OUT[17]),
                      .MU0_MATHB_EFPGA_MAC_OUT_16_(MU0_MATHB_EFPGA_MAC_OUT[16]),
                      .MU0_MATHB_EFPGA_MAC_OUT_15_(MU0_MATHB_EFPGA_MAC_OUT[15]),
                      .MU0_MATHB_EFPGA_MAC_OUT_14_(MU0_MATHB_EFPGA_MAC_OUT[14]),
                      .MU0_MATHB_EFPGA_MAC_OUT_13_(MU0_MATHB_EFPGA_MAC_OUT[13]),
                      .MU0_MATHB_EFPGA_MAC_OUT_12_(MU0_MATHB_EFPGA_MAC_OUT[12]),
                      .MU0_MATHB_EFPGA_MAC_OUT_11_(MU0_MATHB_EFPGA_MAC_OUT[11]),
                      .MU0_MATHB_EFPGA_MAC_OUT_10_(MU0_MATHB_EFPGA_MAC_OUT[10]),
                      .MU0_MATHB_EFPGA_MAC_OUT_9_(MU0_MATHB_EFPGA_MAC_OUT[9]),
                      .MU0_MATHB_EFPGA_MAC_OUT_8_(MU0_MATHB_EFPGA_MAC_OUT[8]),