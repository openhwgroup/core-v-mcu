module a2_bootrom
 #(
 parameter ADDR_WIDTH=32,
 parameter DATA_WIDTH=32
 )
 (
 input logic 		  CLK,
 input logic 		  CEN,
 input logic [ADDR_WIDTH-1:0]  A,
 output logic [DATA_WIDTH-1:0] Q
 );
 logic [31:0] 		  value;
 assign Q = value;
 always @(posedge CLK) begin
  case (A)
  0: value <= 32'h09C0006F;
  1: value <= 32'h0980006F;
  2: value <= 32'h0940006F;
  3: value <= 32'h0900006F;
  4: value <= 32'h08C0006F;
  5: value <= 32'h0880006F;
  6: value <= 32'h0840006F;
  7: value <= 32'h0800006F;
  8: value <= 32'h07C0006F;
  9: value <= 32'h0780006F;
  10: value <= 32'h0740006F;
  11: value <= 32'h0700006F;
  12: value <= 32'h06C0006F;
  13: value <= 32'h0680006F;
  14: value <= 32'h0640006F;
  15: value <= 32'h0600006F;
  16: value <= 32'h05C0006F;
  17: value <= 32'h0580006F;
  18: value <= 32'h0540006F;
  19: value <= 32'h0500006F;
  20: value <= 32'h04C0006F;
  21: value <= 32'h0480006F;
  22: value <= 32'h0440006F;
  23: value <= 32'h0400006F;
  24: value <= 32'h03C0006F;
  25: value <= 32'h0380006F;
  26: value <= 32'h0340006F;
  27: value <= 32'h0300006F;
  28: value <= 32'h02C0006F;
  29: value <= 32'h0280006F;
  30: value <= 32'h0240006F;
  31: value <= 32'h0200006F;
  32: value <= 32'h0080006F;
  33: value <= 32'h0000006F;
  34: value <= 32'h0207E117;
  35: value <= 32'hFE410113;
  36: value <= 32'h4FA0006F;
  37: value <= 32'h00060113;
  38: value <= 32'h00058067;
  39: value <= 32'h30200073;
  40: value <= 32'hCA09832A;
  41: value <= 32'h00058383;
  42: value <= 32'h00730023;
  43: value <= 32'h0305167D;
  44: value <= 32'hFA6D0585;
  45: value <= 32'h11018082;
  46: value <= 32'hE937C84A;
  47: value <= 32'hC4521C07;
  48: value <= 32'hC6990A13;
  49: value <= 32'h4983C64E;
  50: value <= 32'hCC22000A;
  51: value <= 32'hCA26CE06;
  52: value <= 32'h842A4785;
  53: value <= 32'hC6990913;
  54: value <= 32'h06F98563;
  55: value <= 32'h00144783;
  56: value <= 32'h00044703;
  57: value <= 32'h8FD907A2;
  58: value <= 32'h07136729;
  59: value <= 32'h92635077;
  60: value <= 32'h478304E7;
  61: value <= 32'h07130064;
  62: value <= 32'h92630240;
  63: value <= 32'h470308E7;
  64: value <= 32'h47830034;
  65: value <= 32'h45030024;
  66: value <= 32'h07220054;
  67: value <= 32'h47838F5D;
  68: value <= 32'h46030044;
  69: value <= 32'h05620074;
  70: value <= 32'h8FD907C2;
  71: value <= 32'h00840593;
  72: value <= 32'h3FBD8D5D;
  73: value <= 32'h00094703;
  74: value <= 32'h05134785;
  75: value <= 32'h00630310;
  76: value <= 32'h40F204F7;
  77: value <= 32'h44D24462;
  78: value <= 32'h49B24942;
  79: value <= 32'h61054A22;
  80: value <= 32'h84AE8082;
  81: value <= 32'h05C215F9;
  82: value <= 32'h22AD81C1;
  83: value <= 32'hC70394A2;
  84: value <= 32'hC783FFE4;
  85: value <= 32'h0722FFF4;
  86: value <= 32'h07C28FD9;
  87: value <= 32'h8FE383C1;
  88: value <= 32'h4783F6A7;
  89: value <= 32'h96E3000A;
  90: value <= 32'h0513FD37;
  91: value <= 32'h44620300;
  92: value <= 32'h44D240F2;
  93: value <= 32'h49B24942;
  94: value <= 32'h61054A22;
  95: value <= 32'h0713A47D;
  96: value <= 32'h91E30260;
  97: value <= 32'h1537FAE7;
  98: value <= 32'h05131A00;
  99: value <= 32'h2A51A0C5;
  100: value <= 32'h00344703;
  101: value <= 32'h00244783;
  102: value <= 32'h00544503;
  103: value <= 32'h8F5D0722;
  104: value <= 32'h00444783;
  105: value <= 32'h07C20562;
  106: value <= 32'h8D5D8FD9;
  107: value <= 32'h153722CD;
  108: value <= 32'h05131A00;
  109: value <= 32'h22B5A2C5;
  110: value <= 32'h00344783;
  111: value <= 32'h00244703;
  112: value <= 32'h8FD907A2;
  113: value <= 32'h00444703;
  114: value <= 32'h8F5D0742;
  115: value <= 32'h00544783;
  116: value <= 32'h8FD907E2;
  117: value <= 32'hA0019782;
  118: value <= 32'hC6061141;
  119: value <= 32'hC226C422;
  120: value <= 32'h2C35C04A;
  121: value <= 32'hE7B7CD35;
  122: value <= 32'h44051C07;
  123: value <= 32'hC6878423;
  124: value <= 32'h47E5240D;
  125: value <= 32'h00F51E63;
  126: value <= 32'h1C07E7B7;
  127: value <= 32'hC60784A3;
  128: value <= 32'h40B24422;
  129: value <= 32'h49024492;
  130: value <= 32'h02100513;
  131: value <= 32'hAC310141;
  132: value <= 32'h07932409;
  133: value <= 32'h17630200;
  134: value <= 32'hE7B700F5;
  135: value <= 32'h84A31C07;
  136: value <= 32'hBFF9C687;
  137: value <= 32'h079322FD;
  138: value <= 32'h1B630230;
  139: value <= 32'hE4B702F5;
  140: value <= 32'h44011C07;
  141: value <= 32'h92848913;
  142: value <= 32'h2A75A809;
  143: value <= 32'h008907B3;
  144: value <= 32'h04420405;
  145: value <= 32'h00A78023;
  146: value <= 32'h2A6D8041;
  147: value <= 32'h85A2F57D;
  148: value <= 32'h40B24422;
  149: value <= 32'h85134902;
  150: value <= 32'h44929284;
  151: value <= 32'hBDA10141;
  152: value <= 32'h442240B2;
  153: value <= 32'h49024492;
  154: value <= 32'h80820141;
  155: value <= 32'h1C07E737;
  156: value <= 32'h07136585;
  157: value <= 32'h4601A287;
  158: value <= 32'h02158593;
  159: value <= 32'h10000513;
  160: value <= 32'h00861793;
  161: value <= 32'h83C107C2;
  162: value <= 32'h981346A1;
  163: value <= 32'h58130107;
  164: value <= 32'h07864108;
  165: value <= 32'h00085363;
  166: value <= 32'h16FD8FAD;
  167: value <= 32'hF69307C2;
  168: value <= 32'h83C10FF6;
  169: value <= 32'h1023F2FD;
  170: value <= 32'h060500F7;
  171: value <= 32'h19E30709;
  172: value <= 32'h8082FCA6;
  173: value <= 32'hE63767C1;
  174: value <= 32'h86AA1C07;
  175: value <= 32'h85134701;
  176: value <= 32'h0613FFF7;
  177: value <= 32'h4363A286;
  178: value <= 32'h808200B7;
  179: value <= 32'h00E68833;
  180: value <= 32'h00084803;
  181: value <= 32'h00855793;
  182: value <= 32'hC7B30705;
  183: value <= 32'h07860107;
  184: value <= 32'hD80397B2;
  185: value <= 32'h17930007;
  186: value <= 32'h07C20085;
  187: value <= 32'h453383C1;
  188: value <= 32'hBFD100F8;
  189: value <= 32'hC62A1101;
  190: value <= 32'h45850070;
  191: value <= 32'hCE064505;
  192: value <= 32'h40F22DD9;
  193: value <= 32'h80826105;
  194: value <= 32'h45351141;
  195: value <= 32'h37DDC606;
  196: value <= 32'h452940B2;
  197: value <= 32'hBFF90141;
  198: value <= 32'h136347A9;
  199: value <= 32'hB7ED00F5;
  200: value <= 32'h1141BFD1;
  201: value <= 32'hC606C422;
  202: value <= 32'h0503842A;
  203: value <= 32'hE5090004;
  204: value <= 32'h442240B2;
  205: value <= 32'h80820141;
  206: value <= 32'h040537C5;
  207: value <= 32'h5793B7FD;
  208: value <= 32'h11410045;
  209: value <= 32'hC4228BBD;
  210: value <= 32'h842AC606;
  211: value <= 32'h03900713;
  212: value <= 32'h03078513;
  213: value <= 32'h00A75463;
  214: value <= 32'h05778513;
  215: value <= 32'h883D3F75;
  216: value <= 32'h03040513;
  217: value <= 32'h03900793;
  218: value <= 32'h00A7D463;
  219: value <= 32'h05740513;
  220: value <= 32'h40B24422;
  221: value <= 32'hB74D0141;
  222: value <= 32'hC4221141;
  223: value <= 32'h8121842A;
  224: value <= 32'h3F75C606;
  225: value <= 32'h44228522;
  226: value <= 32'h014140B2;
  227: value <= 32'h1141BF4D;
  228: value <= 32'h842AC422;
  229: value <= 32'hC6068141;
  230: value <= 32'h852237C5;
  231: value <= 32'h40B24422;
  232: value <= 32'hBFD90141;
  233: value <= 32'h1A1077B7;
  234: value <= 32'h75134388;
  235: value <= 32'h808207F5;
  236: value <= 32'h1A107737;
  237: value <= 32'h00074783;
  238: value <= 32'h07F57513;
  239: value <= 32'hF807F793;
  240: value <= 32'h00238FC9;
  241: value <= 32'h808200F7;
  242: value <= 32'h1F634785;
  243: value <= 32'h773700F5;
  244: value <= 32'h47831A10;
  245: value <= 32'hE7930047;
  246: value <= 32'h02230017;
  247: value <= 32'h77B700F7;
  248: value <= 32'h43C81A10;
  249: value <= 32'h80828905;
  250: value <= 32'h7737F97D;
  251: value <= 32'h47831A10;
  252: value <= 32'h9BF90047;
  253: value <= 32'h77B7B7DD;
  254: value <= 32'hA5031A10;
  255: value <= 32'h75130847;
  256: value <= 32'h80820FF5;
  257: value <= 32'h1A1077B7;
  258: value <= 32'h0907A503;
  259: value <= 32'h0FF57513;
  260: value <= 32'h77B78082;
  261: value <= 32'h43A81A10;
  262: value <= 32'h0FF57513;
  263: value <= 32'h77B78082;
  264: value <= 32'h43E81A10;
  265: value <= 32'h0FF57513;
  266: value <= 32'h77B78082;
  267: value <= 32'hC7A81A10;
  268: value <= 32'h11418082;
  269: value <= 32'h6485C226;
  270: value <= 32'h40848593;
  271: value <= 32'h4641C422;
  272: value <= 32'h95AA842A;
  273: value <= 32'hC6064501;
  274: value <= 32'h29BD94A2;
  275: value <= 32'h40C4A603;
  276: value <= 32'hCE6347BD;
  277: value <= 32'hCE1100C7;
  278: value <= 32'h85936585;
  279: value <= 32'h95A24185;
  280: value <= 32'h40B24422;
  281: value <= 32'h06124492;
  282: value <= 32'h01414541;
  283: value <= 32'h4641A9B1;
  284: value <= 32'h40B2B7E5;
  285: value <= 32'h44924422;
  286: value <= 32'h80820141;
  287: value <= 32'hD64E7139;
  288: value <= 32'hDA266985;
  289: value <= 32'hD05AD84A;
  290: value <= 32'h8493892A;
  291: value <= 32'h6B094189;
  292: value <= 32'hC86AD256;
  293: value <= 32'hDC22DE06;
  294: value <= 32'hCE5ED452;
  295: value <= 32'hCA66CC62;
  296: value <= 32'h94CAC66E;
  297: value <= 32'h4A813779;
  298: value <= 32'h9B4A99CA;
  299: value <= 32'h01000D37;
  300: value <= 32'h40C9A783;
  301: value <= 32'h02FAE363;
  302: value <= 32'h1A001537;
  303: value <= 32'hA3050513;
  304: value <= 32'hA503358D;
  305: value <= 32'h35E14109;
  306: value <= 32'h1A001537;
  307: value <= 32'hA2C50513;
  308: value <= 32'hA7833D89;
  309: value <= 32'h97824109;
  310: value <= 32'h17B7A001;
  311: value <= 32'h85131A00;
  312: value <= 32'h3581A1C7;
  313: value <= 32'h35658556;
  314: value <= 32'h1A0017B7;
  315: value <= 32'hA3878513;
  316: value <= 32'h40C83D0D;
  317: value <= 32'hE4000BB7;
  318: value <= 32'h3D514C01;
  319: value <= 32'h0044AA03;
  320: value <= 32'h0004AC83;
  321: value <= 32'h0084AD83;
  322: value <= 32'h44D49BD2;
  323: value <= 32'h00DC6563;
  324: value <= 32'h04C10A85;
  325: value <= 32'h2403BF71;
  326: value <= 32'hF563920B;
  327: value <= 32'h8413008D;
  328: value <= 32'h9871003D;
  329: value <= 32'hFB638622;
  330: value <= 32'h85D201AB;
  331: value <= 32'h2E698566;
  332: value <= 32'h9CA29A22;
  333: value <= 32'h408D8DB3;
  334: value <= 32'hBFC10C05;
  335: value <= 32'h856685CA;
  336: value <= 32'h86222661;
  337: value <= 32'h855285CA;
  338: value <= 32'hB7DD3EA1;
  339: value <= 32'h4785C505;
  340: value <= 32'h02F50563;
  341: value <= 32'h17634789;
  342: value <= 32'h07B702F5;
  343: value <= 32'h87931A10;
  344: value <= 32'h43980407;
  345: value <= 32'h000806B7;
  346: value <= 32'hC3988F55;
  347: value <= 32'h9B6D4398;
  348: value <= 32'h8082C398;
  349: value <= 32'h1A1007B7;
  350: value <= 32'h07B7B7ED;
  351: value <= 32'h87931A10;
  352: value <= 32'hB7C50207;
  353: value <= 32'h00002783;
  354: value <= 32'h71799002;
  355: value <= 32'hD6064501;
  356: value <= 32'hD226D422;
  357: value <= 32'hCE4ED04A;
  358: value <= 32'h3F4DCC52;
  359: value <= 32'h377D4505;
  360: value <= 32'h376D4509;
  361: value <= 32'h1C0107B7;
  362: value <= 32'h4505439C;
  363: value <= 32'h1A1047B7;
  364: value <= 32'h0C47A403;
  365: value <= 32'h33FD3D11;
  366: value <= 32'h06200793;
  367: value <= 32'h05638805;
  368: value <= 32'h051300F5;
  369: value <= 32'h33ED0620;
  370: value <= 32'h859365F1;
  371: value <= 32'h45052005;
  372: value <= 32'h1537264D;
  373: value <= 32'h05131A00;
  374: value <= 32'h33A1A405;
  375: value <= 32'h1A001537;
  376: value <= 32'hA4C50513;
  377: value <= 32'h15373B3D;
  378: value <= 32'h05131A00;
  379: value <= 32'h3B15A505;
  380: value <= 32'h1A001537;
  381: value <= 32'hA5C50513;
  382: value <= 32'hC455332D;
  383: value <= 32'h1A001537;
  384: value <= 32'hA7450513;
  385: value <= 32'h25B73B39;
  386: value <= 32'h85930026;
  387: value <= 32'h45015A05;
  388: value <= 32'h45812235;
  389: value <= 32'h22ED4501;
  390: value <= 32'h45014581;
  391: value <= 32'h002824A1;
  392: value <= 32'hE4092A91;
  393: value <= 32'h02E00793;
  394: value <= 32'h00F10423;
  395: value <= 32'h000104A3;
  396: value <= 32'hC537C44D;
  397: value <= 32'h67851C07;
  398: value <= 32'h00050413;
  399: value <= 32'h09336489;
  400: value <= 32'h05130094;
  401: value <= 32'h943E0005;
  402: value <= 32'h92F92023;
  403: value <= 32'h90092E23;
  404: value <= 32'h40042223;
  405: value <= 32'h92092223;
  406: value <= 32'h27833BE9;
  407: value <= 32'h28039209;
  408: value <= 32'hD73740C4;
  409: value <= 32'h88931C07;
  410: value <= 32'h06B3FFF7;
  411: value <= 32'h071340F0;
  412: value <= 32'h46014207;
  413: value <= 32'h1C000537;
  414: value <= 32'h92848493;
  415: value <= 32'h03061A63;
  416: value <= 32'h97AA6789;
  417: value <= 32'hA0236605;
  418: value <= 32'h061392C7;
  419: value <= 32'h962A5196;
  420: value <= 32'h1A0005B7;
  421: value <= 32'h9007AE23;
  422: value <= 32'h9207A223;
  423: value <= 32'h40060613;
  424: value <= 32'h47C58593;
  425: value <= 32'h15373AC5;
  426: value <= 32'h05131A00;
  427: value <= 32'hBF99A785;
  428: value <= 32'hFFC72783;
  429: value <= 32'h00F56963;
  430: value <= 32'h95BE430C;
  431: value <= 32'h00B56963;
  432: value <= 32'h07410605;
  433: value <= 32'h05B3BF65;
  434: value <= 32'hFBE30095;
  435: value <= 32'h430CFEB7;
  436: value <= 32'h97C697AE;
  437: value <= 32'h00D7F533;
  438: value <= 32'h3E49B7E5;
  439: value <= 32'h1A1047B7;
  440: value <= 32'h0DC7A683;
  441: value <= 32'h05134705;
  442: value <= 32'h88630270;
  443: value <= 32'hA78300E6;
  444: value <= 32'h8B890DC7;
  445: value <= 32'h0513C781;
  446: value <= 32'h3B050280;
  447: value <= 32'h1A1047B7;
  448: value <= 32'hDBF84705;
  449: value <= 32'h0007A4B7;
  450: value <= 32'h1A104937;
  451: value <= 32'hEA374985;
  452: value <= 32'h84131C07;
  453: value <= 32'h27831204;
  454: value <= 32'h88630749;
  455: value <= 32'h87B70137;
  456: value <= 32'h87931C00;
  457: value <= 32'h97820807;
  458: value <= 32'h147DA001;
  459: value <= 32'hF4653475;
  460: value <= 32'hC68A4783;
  461: value <= 32'h0028FFF9;
  462: value <= 32'hBFE136ED;
  463: value <= 32'h1A102737;
  464: value <= 32'h47914714;
  465: value <= 32'h00A79533;
  466: value <= 32'hC7148EC9;
  467: value <= 32'h47934714;
  468: value <= 32'h8FF5FFF5;
  469: value <= 32'h431CC71C;
  470: value <= 32'h57B78D5D;
  471: value <= 32'h8793004C;
  472: value <= 32'hD7B3B407;
  473: value <= 32'hC30802B7;
  474: value <= 32'h1C07E737;
  475: value <= 32'h05234501;
  476: value <= 32'h8082C6F7;
  477: value <= 32'h1A102637;
  478: value <= 32'h18864703;
  479: value <= 32'h1C07E6B7;
  480: value <= 32'h18060793;
  481: value <= 32'h04239B3D;
  482: value <= 32'h470318E6;
  483: value <= 32'h9B3D1986;
  484: value <= 32'h18E60C23;
  485: value <= 32'h1A864703;
  486: value <= 32'h04239B3D;
  487: value <= 32'hC6831AE6;
  488: value <= 32'hE737C6A6;
  489: value <= 32'h07131C07;
  490: value <= 32'hC314C287;
  491: value <= 32'h100006B7;
  492: value <= 32'h06B7C354;
  493: value <= 32'h86932007;
  494: value <= 32'hC71409F6;
  495: value <= 32'h704706B7;
  496: value <= 32'hC754068D;
  497: value <= 32'h900006B7;
  498: value <= 32'hCB140685;
  499: value <= 32'h18A62023;
  500: value <= 32'hC3D44691;
  501: value <= 32'h18864683;
  502: value <= 32'h0106E693;
  503: value <= 32'h18D60423;
  504: value <= 32'h4751D398;
  505: value <= 32'h4703D3D8;
  506: value <= 32'h67131A86;
  507: value <= 32'h04230107;
  508: value <= 32'h27371AE6;
  509: value <= 32'h07931A10;
  510: value <= 32'h43DC1807;
  511: value <= 32'h8082FFED;
  512: value <= 32'h003427B7;
  513: value <= 32'h04378793;
  514: value <= 32'h051E953E;
  515: value <= 32'h02854783;
  516: value <= 32'h1C07E737;
  517: value <= 32'hC6A74703;
  518: value <= 32'h04239BBD;
  519: value <= 32'h478302F5;
  520: value <= 32'hE7930285;
  521: value <= 32'h04230407;
  522: value <= 32'hE7B702F5;
  523: value <= 32'h87931C07;
  524: value <= 32'hC398C287;
  525: value <= 32'h10000737;
  526: value <= 32'h07378DD9;
  527: value <= 32'h07132007;
  528: value <= 32'hC7980667;
  529: value <= 32'h90000737;
  530: value <= 32'hD11C0705;
  531: value <= 32'hC7D8C3CC;
  532: value <= 32'hD15C47C1;
  533: value <= 32'h02854783;
  534: value <= 32'h0107E793;
  535: value <= 32'h02F50423;
  536: value <= 32'h80824501;
  537: value <= 32'h003427B7;
  538: value <= 32'h04378793;
  539: value <= 32'h051E953E;
  540: value <= 32'h02854783;
  541: value <= 32'h1C07E737;
  542: value <= 32'hC6A74703;
  543: value <= 32'h04239BBD;
  544: value <= 32'h478302F5;
  545: value <= 32'hE7930285;
  546: value <= 32'h04230407;
  547: value <= 32'hE7B702F5;
  548: value <= 32'h87931C07;
  549: value <= 32'hC398C287;
  550: value <= 32'h10000737;
  551: value <= 32'h07378DD9;
  552: value <= 32'h07132007;
  553: value <= 32'hC7980997;
  554: value <= 32'h90000737;
  555: value <= 32'hD11C0705;
  556: value <= 32'hC7D8C3CC;
  557: value <= 32'hD15C47C1;
  558: value <= 32'h02854783;
  559: value <= 32'h0107E793;
  560: value <= 32'h02F50423;
  561: value <= 32'h80824501;
  562: value <= 32'h1A102837;
  563: value <= 32'h18884703;
  564: value <= 32'h1C07E6B7;
  565: value <= 32'h200708B7;
  566: value <= 32'h04239B3D;
  567: value <= 32'h470318E8;
  568: value <= 32'h03371988;
  569: value <= 32'h0793200F;
  570: value <= 32'h9B3D1808;
  571: value <= 32'h18E80C23;
  572: value <= 32'h1A884703;
  573: value <= 32'h04239B3D;
  574: value <= 32'hC6831AE8;
  575: value <= 32'hE737C6A6;
  576: value <= 32'h07131C07;
  577: value <= 32'hC314C287;
  578: value <= 32'h100006B7;
  579: value <= 32'h8693C354;
  580: value <= 32'hC7140038;
  581: value <= 32'h00855693;
  582: value <= 32'h82C106C2;
  583: value <= 32'h0FF57513;
  584: value <= 32'h0066E6B3;
  585: value <= 32'h01156533;
  586: value <= 32'hCB08C754;
  587: value <= 32'hFFF60693;
  588: value <= 32'h70470537;
  589: value <= 32'hCB548EC9;
  590: value <= 32'h900006B7;
  591: value <= 32'hCF140685;
  592: value <= 32'h18B82023;
  593: value <= 32'h4683C3D0;
  594: value <= 32'hE6931888;
  595: value <= 32'h04230106;
  596: value <= 32'hD39818D8;
  597: value <= 32'hD3D84771;
  598: value <= 32'h1A884703;
  599: value <= 32'h01076713;
  600: value <= 32'h1AE80423;
  601: value <= 32'h1A102737;
  602: value <= 32'h18070793;
  603: value <= 32'hFFED43DC;
  604: value <= 32'h27378082;
  605: value <= 32'h47141A10;
  606: value <= 32'h97B34785;
  607: value <= 32'h8EDD00A7;
  608: value <= 32'h4710C714;
  609: value <= 32'hFFF7C693;
  610: value <= 32'hC7148EF1;
  611: value <= 32'h8FD54314;
  612: value <= 32'h27B7C31C;
  613: value <= 32'h87930034;
  614: value <= 32'h953E0417;
  615: value <= 32'h004C57B7;
  616: value <= 32'hB4078793;
  617: value <= 32'h02B7D7B3;
  618: value <= 32'h07C2051E;
  619: value <= 32'h132383C1;
  620: value <= 32'h515C02F5;
  621: value <= 32'h0067E793;
  622: value <= 32'h515CD15C;
  623: value <= 32'h0107E793;
  624: value <= 32'h515CD15C;
  625: value <= 32'h1007E793;
  626: value <= 32'h515CD15C;
  627: value <= 32'h2007E793;
  628: value <= 32'h4501D15C;
  629: value <= 32'h27B78082;
  630: value <= 32'h87930034;
  631: value <= 32'h953E0417;
  632: value <= 32'h00751793;
  633: value <= 32'h4BD84501;
  634: value <= 32'hCB90EF11;
  635: value <= 32'hC703CBCC;
  636: value <= 32'h67130187;
  637: value <= 32'h8C230107;
  638: value <= 32'h4BD800E7;
  639: value <= 32'h0542E711;
  640: value <= 32'h80828141;
  641: value <= 32'hB7C50505;
  642: value <= 32'hBFC50505;
  643: value <= 32'h4332490A;
  644: value <= 32'h204C4220;
  645: value <= 32'h20504D4A;
  646: value <= 32'h00000000;
  647: value <= 32'h616F4C0A;
  648: value <= 32'h676E6964;
  649: value <= 32'h63655320;
  650: value <= 32'h6E6F6974;
  651: value <= 32'h00000020;
  652: value <= 32'h6D754A0A;
  653: value <= 32'h676E6970;
  654: value <= 32'h206F7420;
  655: value <= 32'h00000000;
  656: value <= 32'h206E614A;
  657: value <= 32'h32203320;
  658: value <= 32'h00323230;
  659: value <= 32'h00002020;
  660: value <= 32'h343A3730;
  661: value <= 32'h32343A30;
  662: value <= 32'h00000000;
  663: value <= 32'h2032410A;
  664: value <= 32'h746F6F42;
  665: value <= 32'h64616F6C;
  666: value <= 32'h42207265;
  667: value <= 32'h73746F6F;
  668: value <= 32'h003D6C65;
  669: value <= 32'h00000031;
  670: value <= 32'h00000030;
  default: value <= 0;
   endcase
  end
endmodule    
