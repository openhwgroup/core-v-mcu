/*****************************************************************
          Vendor       : QuickLogic Corp.
          File Name    : QL_eFPGA_ArcticPro2_32X32_GF_22_top1.vq
          Author       : QuickLogic Corp.

          Description : Verilog Simulation Netlist file
******************************************************************/


module QL_eFPGA_ArcticPro2_32X32_GF_22_Arnold2 (
    input  A2F_B_10_0,
    input  A2F_B_10_1,
    input  A2F_B_10_2,
    input  A2F_B_10_3,
    input  A2F_B_10_4,
    input  A2F_B_10_5,
    input  A2F_B_10_6,
    input  A2F_B_10_7,
    input  A2F_B_11_0,
    input  A2F_B_11_1,
    input  A2F_B_11_2,
    input  A2F_B_11_3,
    input  A2F_B_11_4,
    input  A2F_B_11_5,
    input  A2F_B_12_0,
    input  A2F_B_12_1,
    input  A2F_B_12_2,
    input  A2F_B_12_3,
    input  A2F_B_12_4,
    input  A2F_B_12_5,
    input  A2F_B_12_6,
    input  A2F_B_12_7,
    input  A2F_B_13_0,
    input  A2F_B_13_1,
    input  A2F_B_13_2,
    input  A2F_B_13_3,
    input  A2F_B_13_4,
    input  A2F_B_13_5,
    input  A2F_B_14_0,
    input  A2F_B_14_1,
    input  A2F_B_14_2,
    input  A2F_B_14_3,
    input  A2F_B_14_4,
    input  A2F_B_14_5,
    input  A2F_B_14_6,
    input  A2F_B_14_7,
    input  A2F_B_15_0,
    input  A2F_B_15_1,
    input  A2F_B_15_2,
    input  A2F_B_15_3,
    input  A2F_B_15_4,
    input  A2F_B_15_5,
    input  A2F_B_16_0,
    input  A2F_B_16_1,
    input  A2F_B_16_2,
    input  A2F_B_16_3,
    input  A2F_B_16_4,
    input  A2F_B_16_5,
    input  A2F_B_16_6,
    input  A2F_B_16_7,
    input  A2F_B_17_0,
    input  A2F_B_17_1,
    input  A2F_B_17_2,
    input  A2F_B_17_3,
    input  A2F_B_17_4,
    input  A2F_B_17_5,
    input  A2F_B_18_0,
    input  A2F_B_18_1,
    input  A2F_B_18_2,
    input  A2F_B_18_3,
    input  A2F_B_18_4,
    input  A2F_B_18_5,
    input  A2F_B_18_6,
    input  A2F_B_18_7,
    input  A2F_B_19_0,
    input  A2F_B_19_1,
    input  A2F_B_19_2,
    input  A2F_B_19_3,
    input  A2F_B_19_4,
    input  A2F_B_19_5,
    input  A2F_B_1_0,
    input  A2F_B_1_1,
    input  A2F_B_1_2,
    input  A2F_B_1_3,
    input  A2F_B_1_4,
    input  A2F_B_1_5,
    input  A2F_B_20_0,
    input  A2F_B_20_1,
    input  A2F_B_20_2,
    input  A2F_B_20_3,
    input  A2F_B_20_4,
    input  A2F_B_20_5,
    input  A2F_B_20_6,
    input  A2F_B_20_7,
    input  A2F_B_21_0,
    input  A2F_B_21_1,
    input  A2F_B_21_2,
    input  A2F_B_21_3,
    input  A2F_B_21_4,
    input  A2F_B_21_5,
    input  A2F_B_22_0,
    input  A2F_B_22_1,
    input  A2F_B_22_2,
    input  A2F_B_22_3,
    input  A2F_B_22_4,
    input  A2F_B_22_5,
    input  A2F_B_22_6,
    input  A2F_B_22_7,
    input  A2F_B_23_0,
    input  A2F_B_23_1,
    input  A2F_B_23_2,
    input  A2F_B_23_3,
    input  A2F_B_23_4,
    input  A2F_B_23_5,
    input  A2F_B_24_0,
    input  A2F_B_24_1,
    input  A2F_B_24_2,
    input  A2F_B_24_3,
    input  A2F_B_24_4,
    input  A2F_B_24_5,
    input  A2F_B_24_6,
    input  A2F_B_24_7,
    input  A2F_B_25_0,
    input  A2F_B_25_1,
    input  A2F_B_25_2,
    input  A2F_B_25_3,
    input  A2F_B_25_4,
    input  A2F_B_25_5,
    input  A2F_B_26_0,
    input  A2F_B_26_1,
    input  A2F_B_26_2,
    input  A2F_B_26_3,
    input  A2F_B_26_4,
    input  A2F_B_26_5,
    input  A2F_B_26_6,
    input  A2F_B_26_7,
    input  A2F_B_27_0,
    input  A2F_B_27_1,
    input  A2F_B_27_2,
    input  A2F_B_27_3,
    input  A2F_B_27_4,
    input  A2F_B_27_5,
    input  A2F_B_28_0,
    input  A2F_B_28_1,
    input  A2F_B_28_2,
    input  A2F_B_28_3,
    input  A2F_B_28_4,
    input  A2F_B_28_5,
    input  A2F_B_28_6,
    input  A2F_B_28_7,
    input  A2F_B_29_0,
    input  A2F_B_29_1,
    input  A2F_B_29_2,
    input  A2F_B_29_3,
    input  A2F_B_29_4,
    input  A2F_B_29_5,
    input  A2F_B_2_0,
    input  A2F_B_2_1,
    input  A2F_B_2_2,
    input  A2F_B_2_3,
    input  A2F_B_2_4,
    input  A2F_B_2_5,
    input  A2F_B_2_6,
    input  A2F_B_2_7,
    input  A2F_B_30_0,
    input  A2F_B_30_1,
    input  A2F_B_30_2,
    input  A2F_B_30_3,
    input  A2F_B_30_4,
    input  A2F_B_30_5,
    input  A2F_B_30_6,
    input  A2F_B_30_7,
    input  A2F_B_31_0,
    input  A2F_B_31_1,
    input  A2F_B_31_2,
    input  A2F_B_31_3,
    input  A2F_B_31_4,
    input  A2F_B_31_5,
    input  A2F_B_32_0,
    input  A2F_B_32_1,
    input  A2F_B_32_2,
    input  A2F_B_32_3,
    input  A2F_B_32_4,
    input  A2F_B_32_5,
    input  A2F_B_32_6,
    input  A2F_B_32_7,
    input  A2F_B_3_0,
    input  A2F_B_3_1,
    input  A2F_B_3_2,
    input  A2F_B_3_3,
    input  A2F_B_3_4,
    input  A2F_B_3_5,
    input  A2F_B_4_0,
    input  A2F_B_4_1,
    input  A2F_B_4_2,
    input  A2F_B_4_3,
    input  A2F_B_4_4,
    input  A2F_B_4_5,
    input  A2F_B_4_6,
    input  A2F_B_4_7,
    input  A2F_B_5_0,
    input  A2F_B_5_1,
    input  A2F_B_5_2,
    input  A2F_B_5_3,
    input  A2F_B_5_4,
    input  A2F_B_5_5,
    input  A2F_B_6_0,
    input  A2F_B_6_1,
    input  A2F_B_6_2,
    input  A2F_B_6_3,
    input  A2F_B_6_4,
    input  A2F_B_6_5,
    input  A2F_B_6_6,
    input  A2F_B_6_7,
    input  A2F_B_7_0,
    input  A2F_B_7_1,
    input  A2F_B_7_2,
    input  A2F_B_7_3,
    input  A2F_B_7_4,
    input  A2F_B_7_5,
    input  A2F_B_8_0,
    input  A2F_B_8_1,
    input  A2F_B_8_2,
    input  A2F_B_8_3,
    input  A2F_B_8_4,
    input  A2F_B_8_5,
    input  A2F_B_8_6,
    input  A2F_B_8_7,
    input  A2F_B_9_0,
    input  A2F_B_9_1,
    input  A2F_B_9_2,
    input  A2F_B_9_3,
    input  A2F_B_9_4,
    input  A2F_B_9_5,
    input  A2F_CLK0,
    input  A2F_CLK1,
    input  A2F_CLK2,
    input  A2F_CLK3,
    input  A2F_CLK4,
    input  A2F_CLK5,
    input  A2F_L_10_0,
    input  A2F_L_10_1,
    input  A2F_L_10_2,
    input  A2F_L_10_3,
    input  A2F_L_10_4,
    input  A2F_L_10_5,
    input  A2F_L_10_6,
    input  A2F_L_10_7,
    input  A2F_L_11_0,
    input  A2F_L_11_1,
    input  A2F_L_11_2,
    input  A2F_L_11_3,
    input  A2F_L_11_4,
    input  A2F_L_11_5,
    input  A2F_L_12_0,
    input  A2F_L_12_1,
    input  A2F_L_12_2,
    input  A2F_L_12_3,
    input  A2F_L_12_4,
    input  A2F_L_12_5,
    input  A2F_L_12_6,
    input  A2F_L_12_7,
    input  A2F_L_13_0,
    input  A2F_L_13_1,
    input  A2F_L_13_2,
    input  A2F_L_13_3,
    input  A2F_L_13_4,
    input  A2F_L_13_5,
    input  A2F_L_14_0,
    input  A2F_L_14_1,
    input  A2F_L_14_2,
    input  A2F_L_14_3,
    input  A2F_L_14_4,
    input  A2F_L_14_5,
    input  A2F_L_14_6,
    input  A2F_L_14_7,
    input  A2F_L_15_0,
    input  A2F_L_15_1,
    input  A2F_L_15_2,
    input  A2F_L_15_3,
    input  A2F_L_15_4,
    input  A2F_L_15_5,
    input  A2F_L_16_0,
    input  A2F_L_16_1,
    input  A2F_L_16_2,
    input  A2F_L_16_3,
    input  A2F_L_16_4,
    input  A2F_L_16_5,
    input  A2F_L_16_6,
    input  A2F_L_16_7,
    input  A2F_L_17_0,
    input  A2F_L_17_1,
    input  A2F_L_17_2,
    input  A2F_L_17_3,
    input  A2F_L_17_4,
    input  A2F_L_17_5,
    input  A2F_L_18_0,
    input  A2F_L_18_1,
    input  A2F_L_18_2,
    input  A2F_L_18_3,
    input  A2F_L_18_4,
    input  A2F_L_18_5,
    input  A2F_L_18_6,
    input  A2F_L_18_7,
    input  A2F_L_19_0,
    input  A2F_L_19_1,
    input  A2F_L_19_2,
    input  A2F_L_19_3,
    input  A2F_L_19_4,
    input  A2F_L_19_5,
    input  A2F_L_1_0,
    input  A2F_L_1_1,
    input  A2F_L_1_2,
    input  A2F_L_1_3,
    input  A2F_L_1_4,
    input  A2F_L_1_5,
    input  A2F_L_20_0,
    input  A2F_L_20_1,
    input  A2F_L_20_2,
    input  A2F_L_20_3,
    input  A2F_L_20_4,
    input  A2F_L_20_5,
    input  A2F_L_20_6,
    input  A2F_L_20_7,
    input  A2F_L_21_0,
    input  A2F_L_21_1,
    input  A2F_L_21_2,
    input  A2F_L_21_3,
    input  A2F_L_21_4,
    input  A2F_L_21_5,
    input  A2F_L_22_0,
    input  A2F_L_22_1,
    input  A2F_L_22_2,
    input  A2F_L_22_3,
    input  A2F_L_22_4,
    input  A2F_L_22_5,
    input  A2F_L_22_6,
    input  A2F_L_22_7,
    input  A2F_L_23_0,
    input  A2F_L_23_1,
    input  A2F_L_23_2,
    input  A2F_L_23_3,
    input  A2F_L_23_4,
    input  A2F_L_23_5,
    input  A2F_L_24_0,
    input  A2F_L_24_1,
    input  A2F_L_24_2,
    input  A2F_L_24_3,
    input  A2F_L_24_4,
    input  A2F_L_24_5,
    input  A2F_L_24_6,
    input  A2F_L_24_7,
    input  A2F_L_25_0,
    input  A2F_L_25_1,
    input  A2F_L_25_2,
    input  A2F_L_25_3,
    input  A2F_L_25_4,
    input  A2F_L_25_5,
    input  A2F_L_26_0,
    input  A2F_L_26_1,
    input  A2F_L_26_2,
    input  A2F_L_26_3,
    input  A2F_L_26_4,
    input  A2F_L_26_5,
    input  A2F_L_26_6,
    input  A2F_L_26_7,
    input  A2F_L_27_0,
    input  A2F_L_27_1,
    input  A2F_L_27_2,
    input  A2F_L_27_3,
    input  A2F_L_27_4,
    input  A2F_L_27_5,
    input  A2F_L_28_0,
    input  A2F_L_28_1,
    input  A2F_L_28_2,
    input  A2F_L_28_3,
    input  A2F_L_28_4,
    input  A2F_L_28_5,
    input  A2F_L_28_6,
    input  A2F_L_28_7,
    input  A2F_L_29_0,
    input  A2F_L_29_1,
    input  A2F_L_29_2,
    input  A2F_L_29_3,
    input  A2F_L_29_4,
    input  A2F_L_29_5,
    input  A2F_L_2_0,
    input  A2F_L_2_1,
    input  A2F_L_2_2,
    input  A2F_L_2_3,
    input  A2F_L_2_4,
    input  A2F_L_2_5,
    input  A2F_L_2_6,
    input  A2F_L_2_7,
    input  A2F_L_30_0,
    input  A2F_L_30_1,
    input  A2F_L_30_2,
    input  A2F_L_30_3,
    input  A2F_L_30_4,
    input  A2F_L_30_5,
    input  A2F_L_30_6,
    input  A2F_L_30_7,
    input  A2F_L_31_0,
    input  A2F_L_31_1,
    input  A2F_L_31_2,
    input  A2F_L_31_3,
    input  A2F_L_31_4,
    input  A2F_L_31_5,
    input  A2F_L_32_0,
    input  A2F_L_32_1,
    input  A2F_L_32_2,
    input  A2F_L_32_3,
    input  A2F_L_32_4,
    input  A2F_L_32_5,
    input  A2F_L_32_6,
    input  A2F_L_32_7,
    input  A2F_L_3_0,
    input  A2F_L_3_1,
    input  A2F_L_3_2,
    input  A2F_L_3_3,
    input  A2F_L_3_4,
    input  A2F_L_3_5,
    input  A2F_L_4_0,
    input  A2F_L_4_1,
    input  A2F_L_4_2,
    input  A2F_L_4_3,
    input  A2F_L_4_4,
    input  A2F_L_4_5,
    input  A2F_L_4_6,
    input  A2F_L_4_7,
    input  A2F_L_5_0,
    input  A2F_L_5_1,
    input  A2F_L_5_2,
    input  A2F_L_5_3,
    input  A2F_L_5_4,
    input  A2F_L_5_5,
    input  A2F_L_6_0,
    input  A2F_L_6_1,
    input  A2F_L_6_2,
    input  A2F_L_6_3,
    input  A2F_L_6_4,
    input  A2F_L_6_5,
    input  A2F_L_6_6,
    input  A2F_L_6_7,
    input  A2F_L_7_0,
    input  A2F_L_7_1,
    input  A2F_L_7_2,
    input  A2F_L_7_3,
    input  A2F_L_7_4,
    input  A2F_L_7_5,
    input  A2F_L_8_0,
    input  A2F_L_8_1,
    input  A2F_L_8_2,
    input  A2F_L_8_3,
    input  A2F_L_8_4,
    input  A2F_L_8_5,
    input  A2F_L_8_6,
    input  A2F_L_8_7,
    input  A2F_L_9_0,
    input  A2F_L_9_1,
    input  A2F_L_9_2,
    input  A2F_L_9_3,
    input  A2F_L_9_4,
    input  A2F_L_9_5,
    input  A2F_R_10_0,
    input  A2F_R_10_1,
    input  A2F_R_10_2,
    input  A2F_R_10_3,
    input  A2F_R_10_4,
    input  A2F_R_10_5,
    input  A2F_R_10_6,
    input  A2F_R_10_7,
    input  A2F_R_11_0,
    input  A2F_R_11_1,
    input  A2F_R_11_2,
    input  A2F_R_11_3,
    input  A2F_R_11_4,
    input  A2F_R_11_5,
    input  A2F_R_12_0,
    input  A2F_R_12_1,
    input  A2F_R_12_2,
    input  A2F_R_12_3,
    input  A2F_R_12_4,
    input  A2F_R_12_5,
    input  A2F_R_12_6,
    input  A2F_R_12_7,
    input  A2F_R_13_0,
    input  A2F_R_13_1,
    input  A2F_R_13_2,
    input  A2F_R_13_3,
    input  A2F_R_13_4,
    input  A2F_R_13_5,
    input  A2F_R_14_0,
    input  A2F_R_14_1,
    input  A2F_R_14_2,
    input  A2F_R_14_3,
    input  A2F_R_14_4,
    input  A2F_R_14_5,
    input  A2F_R_14_6,
    input  A2F_R_14_7,
    input  A2F_R_15_0,
    input  A2F_R_15_1,
    input  A2F_R_15_2,
    input  A2F_R_15_3,
    input  A2F_R_15_4,
    input  A2F_R_15_5,
    input  A2F_R_16_0,
    input  A2F_R_16_1,
    input  A2F_R_16_2,
    input  A2F_R_16_3,
    input  A2F_R_16_4,
    input  A2F_R_16_5,
    input  A2F_R_16_6,
    input  A2F_R_16_7,
    input  A2F_R_17_0,
    input  A2F_R_17_1,
    input  A2F_R_17_2,
    input  A2F_R_17_3,
    input  A2F_R_17_4,
    input  A2F_R_17_5,
    input  A2F_R_18_0,
    input  A2F_R_18_1,
    input  A2F_R_18_2,
    input  A2F_R_18_3,
    input  A2F_R_18_4,
    input  A2F_R_18_5,
    input  A2F_R_18_6,
    input  A2F_R_18_7,
    input  A2F_R_19_0,
    input  A2F_R_19_1,
    input  A2F_R_19_2,
    input  A2F_R_19_3,
    input  A2F_R_19_4,
    input  A2F_R_19_5,
    input  A2F_R_1_0,
    input  A2F_R_1_1,
    input  A2F_R_1_2,
    input  A2F_R_1_3,
    input  A2F_R_1_4,
    input  A2F_R_1_5,
    input  A2F_R_20_0,
    input  A2F_R_20_1,
    input  A2F_R_20_2,
    input  A2F_R_20_3,
    input  A2F_R_20_4,
    input  A2F_R_20_5,
    input  A2F_R_20_6,
    input  A2F_R_20_7,
    input  A2F_R_21_0,
    input  A2F_R_21_1,
    input  A2F_R_21_2,
    input  A2F_R_21_3,
    input  A2F_R_21_4,
    input  A2F_R_21_5,
    input  A2F_R_22_0,
    input  A2F_R_22_1,
    input  A2F_R_22_2,
    input  A2F_R_22_3,
    input  A2F_R_22_4,
    input  A2F_R_22_5,
    input  A2F_R_22_6,
    input  A2F_R_22_7,
    input  A2F_R_23_0,
    input  A2F_R_23_1,
    input  A2F_R_23_2,
    input  A2F_R_23_3,
    input  A2F_R_23_4,
    input  A2F_R_23_5,
    input  A2F_R_24_0,
    input  A2F_R_24_1,
    input  A2F_R_24_2,
    input  A2F_R_24_3,
    input  A2F_R_24_4,
    input  A2F_R_24_5,
    input  A2F_R_24_6,
    input  A2F_R_24_7,
    input  A2F_R_25_0,
    input  A2F_R_25_1,
    input  A2F_R_25_2,
    input  A2F_R_25_3,
    input  A2F_R_25_4,
    input  A2F_R_25_5,
    input  A2F_R_26_0,
    input  A2F_R_26_1,
    input  A2F_R_26_2,
    input  A2F_R_26_3,
    input  A2F_R_26_4,
    input  A2F_R_26_5,
    input  A2F_R_26_6,
    input  A2F_R_26_7,
    input  A2F_R_27_0,
    input  A2F_R_27_1,
    input  A2F_R_27_2,
    input  A2F_R_27_3,
    input  A2F_R_27_4,
    input  A2F_R_27_5,
    input  A2F_R_28_0,
    input  A2F_R_28_1,
    input  A2F_R_28_2,
    input  A2F_R_28_3,
    input  A2F_R_28_4,
    input  A2F_R_28_5,
    input  A2F_R_28_6,
    input  A2F_R_28_7,
    input  A2F_R_29_0,
    input  A2F_R_29_1,
    input  A2F_R_29_2,
    input  A2F_R_29_3,
    input  A2F_R_29_4,
    input  A2F_R_29_5,
    input  A2F_R_2_0,
    input  A2F_R_2_1,
    input  A2F_R_2_2,
    input  A2F_R_2_3,
    input  A2F_R_2_4,
    input  A2F_R_2_5,
    input  A2F_R_2_6,
    input  A2F_R_2_7,
    input  A2F_R_30_0,
    input  A2F_R_30_1,
    input  A2F_R_30_2,
    input  A2F_R_30_3,
    input  A2F_R_30_4,
    input  A2F_R_30_5,
    input  A2F_R_30_6,
    input  A2F_R_30_7,
    input  A2F_R_31_0,
    input  A2F_R_31_1,
    input  A2F_R_31_2,
    input  A2F_R_31_3,
    input  A2F_R_31_4,
    input  A2F_R_31_5,
    input  A2F_R_32_0,
    input  A2F_R_32_1,
    input  A2F_R_32_2,
    input  A2F_R_32_3,
    input  A2F_R_32_4,
    input  A2F_R_32_5,
    input  A2F_R_32_6,
    input  A2F_R_32_7,
    input  A2F_R_3_0,
    input  A2F_R_3_1,
    input  A2F_R_3_2,
    input  A2F_R_3_3,
    input  A2F_R_3_4,
    input  A2F_R_3_5,
    input  A2F_R_4_0,
    input  A2F_R_4_1,
    input  A2F_R_4_2,
    input  A2F_R_4_3,
    input  A2F_R_4_4,
    input  A2F_R_4_5,
    input  A2F_R_4_6,
    input  A2F_R_4_7,
    input  A2F_R_5_0,
    input  A2F_R_5_1,
    input  A2F_R_5_2,
    input  A2F_R_5_3,
    input  A2F_R_5_4,
    input  A2F_R_5_5,
    input  A2F_R_6_0,
    input  A2F_R_6_1,
    input  A2F_R_6_2,
    input  A2F_R_6_3,
    input  A2F_R_6_4,
    input  A2F_R_6_5,
    input  A2F_R_6_6,
    input  A2F_R_6_7,
    input  A2F_R_7_0,
    input  A2F_R_7_1,
    input  A2F_R_7_2,
    input  A2F_R_7_3,
    input  A2F_R_7_4,
    input  A2F_R_7_5,
    input  A2F_R_8_0,
    input  A2F_R_8_1,
    input  A2F_R_8_2,
    input  A2F_R_8_3,
    input  A2F_R_8_4,
    input  A2F_R_8_5,
    input  A2F_R_8_6,
    input  A2F_R_8_7,
    input  A2F_R_9_0,
    input  A2F_R_9_1,
    input  A2F_R_9_2,
    input  A2F_R_9_3,
    input  A2F_R_9_4,
    input  A2F_R_9_5,
    input  A2F_T_10_0,
    input  A2F_T_10_1,
    input  A2F_T_10_2,
    input  A2F_T_10_3,
    input  A2F_T_10_4,
    input  A2F_T_10_5,
    input  A2F_T_10_6,
    input  A2F_T_10_7,
    input  A2F_T_11_0,
    input  A2F_T_11_1,
    input  A2F_T_11_2,
    input  A2F_T_11_3,
    input  A2F_T_11_4,
    input  A2F_T_11_5,
    input  A2F_T_12_0,
    input  A2F_T_12_1,
    input  A2F_T_12_2,
    input  A2F_T_12_3,
    input  A2F_T_12_4,
    input  A2F_T_12_5,
    input  A2F_T_12_6,
    input  A2F_T_12_7,
    input  A2F_T_13_0,
    input  A2F_T_13_1,
    input  A2F_T_13_2,
    input  A2F_T_13_3,
    input  A2F_T_13_4,
    input  A2F_T_13_5,
    input  A2F_T_14_0,
    input  A2F_T_14_1,
    input  A2F_T_14_2,
    input  A2F_T_14_3,
    input  A2F_T_14_4,
    input  A2F_T_14_5,
    input  A2F_T_14_6,
    input  A2F_T_14_7,
    input  A2F_T_15_0,
    input  A2F_T_15_1,
    input  A2F_T_15_2,
    input  A2F_T_15_3,
    input  A2F_T_15_4,
    input  A2F_T_15_5,
    input  A2F_T_16_0,
    input  A2F_T_16_1,
    input  A2F_T_16_2,
    input  A2F_T_16_3,
    input  A2F_T_16_4,
    input  A2F_T_16_5,
    input  A2F_T_16_6,
    input  A2F_T_16_7,
    input  A2F_T_17_0,
    input  A2F_T_17_1,
    input  A2F_T_17_2,
    input  A2F_T_17_3,
    input  A2F_T_17_4,
    input  A2F_T_17_5,
    input  A2F_T_18_0,
    input  A2F_T_18_1,
    input  A2F_T_18_2,
    input  A2F_T_18_3,
    input  A2F_T_18_4,
    input  A2F_T_18_5,
    input  A2F_T_18_6,
    input  A2F_T_18_7,
    input  A2F_T_19_0,
    input  A2F_T_19_1,
    input  A2F_T_19_2,
    input  A2F_T_19_3,
    input  A2F_T_19_4,
    input  A2F_T_19_5,
    input  A2F_T_1_0,
    input  A2F_T_1_1,
    input  A2F_T_1_2,
    input  A2F_T_1_3,
    input  A2F_T_1_4,
    input  A2F_T_1_5,
    input  A2F_T_20_0,
    input  A2F_T_20_1,
    input  A2F_T_20_2,
    input  A2F_T_20_3,
    input  A2F_T_20_4,
    input  A2F_T_20_5,
    input  A2F_T_20_6,
    input  A2F_T_20_7,
    input  A2F_T_21_0,
    input  A2F_T_21_1,
    input  A2F_T_21_2,
    input  A2F_T_21_3,
    input  A2F_T_21_4,
    input  A2F_T_21_5,
    input  A2F_T_22_0,
    input  A2F_T_22_1,
    input  A2F_T_22_2,
    input  A2F_T_22_3,
    input  A2F_T_22_4,
    input  A2F_T_22_5,
    input  A2F_T_22_6,
    input  A2F_T_22_7,
    input  A2F_T_23_0,
    input  A2F_T_23_1,
    input  A2F_T_23_2,
    input  A2F_T_23_3,
    input  A2F_T_23_4,
    input  A2F_T_23_5,
    input  A2F_T_24_0,
    input  A2F_T_24_1,
    input  A2F_T_24_2,
    input  A2F_T_24_3,
    input  A2F_T_24_4,
    input  A2F_T_24_5,
    input  A2F_T_24_6,
    input  A2F_T_24_7,
    input  A2F_T_25_0,
    input  A2F_T_25_1,
    input  A2F_T_25_2,
    input  A2F_T_25_3,
    input  A2F_T_25_4,
    input  A2F_T_25_5,
    input  A2F_T_26_0,
    input  A2F_T_26_1,
    input  A2F_T_26_2,
    input  A2F_T_26_3,
    input  A2F_T_26_4,
    input  A2F_T_26_5,
    input  A2F_T_26_6,
    input  A2F_T_26_7,
    input  A2F_T_27_0,
    input  A2F_T_27_1,
    input  A2F_T_27_2,
    input  A2F_T_27_3,
    input  A2F_T_27_4,
    input  A2F_T_27_5,
    input  A2F_T_28_0,
    input  A2F_T_28_1,
    input  A2F_T_28_2,
    input  A2F_T_28_3,
    input  A2F_T_28_4,
    input  A2F_T_28_5,
    input  A2F_T_28_6,
    input  A2F_T_28_7,
    input  A2F_T_29_0,
    input  A2F_T_29_1,
    input  A2F_T_29_2,
    input  A2F_T_29_3,
    input  A2F_T_29_4,
    input  A2F_T_29_5,
    input  A2F_T_2_0,
    input  A2F_T_2_1,
    input  A2F_T_2_2,
    input  A2F_T_2_3,
    input  A2F_T_2_4,
    input  A2F_T_2_5,
    input  A2F_T_2_6,
    input  A2F_T_2_7,
    input  A2F_T_30_0,
    input  A2F_T_30_1,
    input  A2F_T_30_2,
    input  A2F_T_30_3,
    input  A2F_T_30_4,
    input  A2F_T_30_5,
    input  A2F_T_30_6,
    input  A2F_T_30_7,
    input  A2F_T_31_0,
    input  A2F_T_31_1,
    input  A2F_T_31_2,
    input  A2F_T_31_3,
    input  A2F_T_31_4,
    input  A2F_T_31_5,
    input  A2F_T_32_0,
    input  A2F_T_32_1,
    input  A2F_T_32_2,
    input  A2F_T_32_3,
    input  A2F_T_32_4,
    input  A2F_T_32_5,
    input  A2F_T_32_6,
    input  A2F_T_32_7,
    input  A2F_T_3_0,
    input  A2F_T_3_1,
    input  A2F_T_3_2,
    input  A2F_T_3_3,
    input  A2F_T_3_4,
    input  A2F_T_3_5,
    input  A2F_T_4_0,
    input  A2F_T_4_1,
    input  A2F_T_4_2,
    input  A2F_T_4_3,
    input  A2F_T_4_4,
    input  A2F_T_4_5,
    input  A2F_T_4_6,
    input  A2F_T_4_7,
    input  A2F_T_5_0,
    input  A2F_T_5_1,
    input  A2F_T_5_2,
    input  A2F_T_5_3,
    input  A2F_T_5_4,
    input  A2F_T_5_5,
    input  A2F_T_6_0,
    input  A2F_T_6_1,
    input  A2F_T_6_2,
    input  A2F_T_6_3,
    input  A2F_T_6_4,
    input  A2F_T_6_5,
    input  A2F_T_6_6,
    input  A2F_T_6_7,
    input  A2F_T_7_0,
    input  A2F_T_7_1,
    input  A2F_T_7_2,
    input  A2F_T_7_3,
    input  A2F_T_7_4,
    input  A2F_T_7_5,
    input  A2F_T_8_0,
    input  A2F_T_8_1,
    input  A2F_T_8_2,
    input  A2F_T_8_3,
    input  A2F_T_8_4,
    input  A2F_T_8_5,
    input  A2F_T_8_6,
    input  A2F_T_8_7,
    input  A2F_T_9_0,
    input  A2F_T_9_1,
    input  A2F_T_9_2,
    input  A2F_T_9_3,
    input  A2F_T_9_4,
    input  A2F_T_9_5,
    input  A2Freg_B_11_0,
    input  A2Freg_B_13_0,
    input  A2Freg_B_15_0,
    input  A2Freg_B_17_0,
    input  A2Freg_B_19_0,
    input  A2Freg_B_1_0,
    input  A2Freg_B_21_0,
    input  A2Freg_B_23_0,
    input  A2Freg_B_25_0,
    input  A2Freg_B_27_0,
    input  A2Freg_B_29_0,
    input  A2Freg_B_31_0,
    input  A2Freg_B_3_0,
    input  A2Freg_B_5_0,
    input  A2Freg_B_7_0,
    input  A2Freg_B_9_0,
    input  A2Freg_L_11_0,
    input  A2Freg_L_13_0,
    input  A2Freg_L_15_0,
    input  A2Freg_L_17_0,
    input  A2Freg_L_19_0,
    input  A2Freg_L_1_0,
    input  A2Freg_L_21_0,
    input  A2Freg_L_23_0,
    input  A2Freg_L_25_0,
    input  A2Freg_L_27_0,
    input  A2Freg_L_29_0,
    input  A2Freg_L_31_0,
    input  A2Freg_L_3_0,
    input  A2Freg_L_5_0,
    input  A2Freg_L_7_0,
    input  A2Freg_L_9_0,
    input  A2Freg_R_11_0,
    input  A2Freg_R_13_0,
    input  A2Freg_R_15_0,
    input  A2Freg_R_17_0,
    input  A2Freg_R_19_0,
    input  A2Freg_R_1_0,
    input  A2Freg_R_21_0,
    input  A2Freg_R_23_0,
    input  A2Freg_R_25_0,
    input  A2Freg_R_27_0,
    input  A2Freg_R_29_0,
    input  A2Freg_R_31_0,
    input  A2Freg_R_3_0,
    input  A2Freg_R_5_0,
    input  A2Freg_R_7_0,
    input  A2Freg_R_9_0,
    input  A2Freg_T_11_0,
    input  A2Freg_T_13_0,
    input  A2Freg_T_15_0,
    input  A2Freg_T_17_0,
    input  A2Freg_T_19_0,
    input  A2Freg_T_1_0,
    input  A2Freg_T_21_0,
    input  A2Freg_T_23_0,
    input  A2Freg_T_25_0,
    input  A2Freg_T_27_0,
    input  A2Freg_T_29_0,
    input  A2Freg_T_31_0,
    input  A2Freg_T_3_0,
    input  A2Freg_T_5_0,
    input  A2Freg_T_7_0,
    input  A2Freg_T_9_0,
    output F2A_B_10_0,
    output F2A_B_10_1,
    output F2A_B_10_10,
    output F2A_B_10_11,
    output F2A_B_10_12,
    output F2A_B_10_13,
    output F2A_B_10_14,
    output F2A_B_10_15,
    output F2A_B_10_16,
    output F2A_B_10_17,
    output F2A_B_10_2,
    output F2A_B_10_3,
    output F2A_B_10_4,
    output F2A_B_10_5,
    output F2A_B_10_6,
    output F2A_B_10_7,
    output F2A_B_10_8,
    output F2A_B_10_9,
    output F2A_B_11_0,
    output F2A_B_11_1,
    output F2A_B_11_10,
    output F2A_B_11_11,
    output F2A_B_11_2,
    output F2A_B_11_3,
    output F2A_B_11_4,
    output F2A_B_11_5,
    output F2A_B_11_6,
    output F2A_B_11_7,
    output F2A_B_11_8,
    output F2A_B_11_9,
    output F2A_B_12_0,
    output F2A_B_12_1,
    output F2A_B_12_10,
    output F2A_B_12_11,
    output F2A_B_12_12,
    output F2A_B_12_13,
    output F2A_B_12_14,
    output F2A_B_12_15,
    output F2A_B_12_16,
    output F2A_B_12_17,
    output F2A_B_12_2,
    output F2A_B_12_3,
    output F2A_B_12_4,
    output F2A_B_12_5,
    output F2A_B_12_6,
    output F2A_B_12_7,
    output F2A_B_12_8,
    output F2A_B_12_9,
    output F2A_B_13_0,
    output F2A_B_13_1,
    output F2A_B_13_10,
    output F2A_B_13_11,
    output F2A_B_13_2,
    output F2A_B_13_3,
    output F2A_B_13_4,
    output F2A_B_13_5,
    output F2A_B_13_6,
    output F2A_B_13_7,
    output F2A_B_13_8,
    output F2A_B_13_9,
    output F2A_B_14_0,
    output F2A_B_14_1,
    output F2A_B_14_10,
    output F2A_B_14_11,
    output F2A_B_14_12,
    output F2A_B_14_13,
    output F2A_B_14_14,
    output F2A_B_14_15,
    output F2A_B_14_16,
    output F2A_B_14_17,
    output F2A_B_14_2,
    output F2A_B_14_3,
    output F2A_B_14_4,
    output F2A_B_14_5,
    output F2A_B_14_6,
    output F2A_B_14_7,
    output F2A_B_14_8,
    output F2A_B_14_9,
    output F2A_B_15_0,
    output F2A_B_15_1,
    output F2A_B_15_10,
    output F2A_B_15_11,
    output F2A_B_15_2,
    output F2A_B_15_3,
    output F2A_B_15_4,
    output F2A_B_15_5,
    output F2A_B_15_6,
    output F2A_B_15_7,
    output F2A_B_15_8,
    output F2A_B_15_9,
    output F2A_B_16_0,
    output F2A_B_16_1,
    output F2A_B_16_10,
    output F2A_B_16_11,
    output F2A_B_16_12,
    output F2A_B_16_13,
    output F2A_B_16_17,
    output F2A_B_16_2,
    output F2A_B_16_3,
    output F2A_B_16_4,
    output F2A_B_16_5,
    output F2A_B_16_6,
    output F2A_B_16_7,
    output F2A_B_16_8,
    output F2A_B_16_9,
    output F2A_B_17_0,
    output F2A_B_17_1,
    output F2A_B_17_10,
    output F2A_B_17_11,
    output F2A_B_17_2,
    output F2A_B_17_3,
    output F2A_B_17_4,
    output F2A_B_17_5,
    output F2A_B_17_6,
    output F2A_B_17_7,
    output F2A_B_17_8,
    output F2A_B_17_9,
    output F2A_B_18_0,
    output F2A_B_18_1,
    output F2A_B_18_10,
    output F2A_B_18_11,
    output F2A_B_18_12,
    output F2A_B_18_13,
    output F2A_B_18_14,
    output F2A_B_18_15,
    output F2A_B_18_16,
    output F2A_B_18_17,
    output F2A_B_18_2,
    output F2A_B_18_3,
    output F2A_B_18_4,
    output F2A_B_18_5,
    output F2A_B_18_6,
    output F2A_B_18_7,
    output F2A_B_18_8,
    output F2A_B_18_9,
    output F2A_B_19_0,
    output F2A_B_19_1,
    output F2A_B_19_10,
    output F2A_B_19_11,
    output F2A_B_19_2,
    output F2A_B_19_3,
    output F2A_B_19_4,
    output F2A_B_19_5,
    output F2A_B_19_6,
    output F2A_B_19_7,
    output F2A_B_19_8,
    output F2A_B_19_9,
    output F2A_B_1_0,
    output F2A_B_1_1,
    output F2A_B_1_10,
    output F2A_B_1_11,
    output F2A_B_1_2,
    output F2A_B_1_3,
    output F2A_B_1_4,
    output F2A_B_1_5,
    output F2A_B_1_6,
    output F2A_B_1_7,
    output F2A_B_1_8,
    output F2A_B_1_9,
    output F2A_B_20_0,
    output F2A_B_20_1,
    output F2A_B_20_10,
    output F2A_B_20_11,
    output F2A_B_20_12,
    output F2A_B_20_13,
    output F2A_B_20_14,
    output F2A_B_20_15,
    output F2A_B_20_16,
    output F2A_B_20_17,
    output F2A_B_20_2,
    output F2A_B_20_3,
    output F2A_B_20_4,
    output F2A_B_20_5,
    output F2A_B_20_6,
    output F2A_B_20_7,
    output F2A_B_20_8,
    output F2A_B_20_9,
    output F2A_B_21_0,
    output F2A_B_21_1,
    output F2A_B_21_10,
    output F2A_B_21_11,
    output F2A_B_21_2,
    output F2A_B_21_3,
    output F2A_B_21_4,
    output F2A_B_21_5,
    output F2A_B_21_6,
    output F2A_B_21_7,
    output F2A_B_21_8,
    output F2A_B_21_9,
    output F2A_B_22_0,
    output F2A_B_22_1,
    output F2A_B_22_10,
    output F2A_B_22_11,
    output F2A_B_22_12,
    output F2A_B_22_13,
    output F2A_B_22_14,
    output F2A_B_22_15,
    output F2A_B_22_16,
    output F2A_B_22_17,
    output F2A_B_22_2,
    output F2A_B_22_3,
    output F2A_B_22_4,
    output F2A_B_22_5,
    output F2A_B_22_6,
    output F2A_B_22_7,
    output F2A_B_22_8,
    output F2A_B_22_9,
    output F2A_B_23_0,
    output F2A_B_23_1,
    output F2A_B_23_10,
    output F2A_B_23_11,
    output F2A_B_23_2,
    output F2A_B_23_3,
    output F2A_B_23_4,
    output F2A_B_23_5,
    output F2A_B_23_6,
    output F2A_B_23_7,
    output F2A_B_23_8,
    output F2A_B_23_9,
    output F2A_B_24_0,
    output F2A_B_24_1,
    output F2A_B_24_10,
    output F2A_B_24_11,
    output F2A_B_24_12,
    output F2A_B_24_13,
    output F2A_B_24_14,
    output F2A_B_24_15,
    output F2A_B_24_16,
    output F2A_B_24_17,
    output F2A_B_24_2,
    output F2A_B_24_3,
    output F2A_B_24_4,
    output F2A_B_24_5,
    output F2A_B_24_6,
    output F2A_B_24_7,
    output F2A_B_24_8,
    output F2A_B_24_9,
    output F2A_B_25_0,
    output F2A_B_25_1,
    output F2A_B_25_10,
    output F2A_B_25_11,
    output F2A_B_25_2,
    output F2A_B_25_3,
    output F2A_B_25_4,
    output F2A_B_25_5,
    output F2A_B_25_6,
    output F2A_B_25_7,
    output F2A_B_25_8,
    output F2A_B_25_9,
    output F2A_B_26_0,
    output F2A_B_26_1,
    output F2A_B_26_10,
    output F2A_B_26_11,
    output F2A_B_26_12,
    output F2A_B_26_13,
    output F2A_B_26_14,
    output F2A_B_26_15,
    output F2A_B_26_16,
    output F2A_B_26_17,
    output F2A_B_26_2,
    output F2A_B_26_3,
    output F2A_B_26_4,
    output F2A_B_26_5,
    output F2A_B_26_6,
    output F2A_B_26_7,
    output F2A_B_26_8,
    output F2A_B_26_9,
    output F2A_B_27_0,
    output F2A_B_27_1,
    output F2A_B_27_10,
    output F2A_B_27_11,
    output F2A_B_27_2,
    output F2A_B_27_3,
    output F2A_B_27_4,
    output F2A_B_27_5,
    output F2A_B_27_6,
    output F2A_B_27_7,
    output F2A_B_27_8,
    output F2A_B_27_9,
    output F2A_B_28_0,
    output F2A_B_28_1,
    output F2A_B_28_10,
    output F2A_B_28_11,
    output F2A_B_28_12,
    output F2A_B_28_13,
    output F2A_B_28_14,
    output F2A_B_28_15,
    output F2A_B_28_16,
    output F2A_B_28_17,
    output F2A_B_28_2,
    output F2A_B_28_3,
    output F2A_B_28_4,
    output F2A_B_28_5,
    output F2A_B_28_6,
    output F2A_B_28_7,
    output F2A_B_28_8,
    output F2A_B_28_9,
    output F2A_B_29_0,
    output F2A_B_29_1,
    output F2A_B_29_10,
    output F2A_B_29_11,
    output F2A_B_29_2,
    output F2A_B_29_3,
    output F2A_B_29_4,
    output F2A_B_29_5,
    output F2A_B_29_6,
    output F2A_B_29_7,
    output F2A_B_29_8,
    output F2A_B_29_9,
    output F2A_B_2_0,
    output F2A_B_2_1,
    output F2A_B_2_10,
    output F2A_B_2_11,
    output F2A_B_2_12,
    output F2A_B_2_13,
    output F2A_B_2_14,
    output F2A_B_2_15,
    output F2A_B_2_16,
    output F2A_B_2_17,
    output F2A_B_2_2,
    output F2A_B_2_3,
    output F2A_B_2_4,
    output F2A_B_2_5,
    output F2A_B_2_6,
    output F2A_B_2_7,
    output F2A_B_2_8,
    output F2A_B_2_9,
    output F2A_B_30_0,
    output F2A_B_30_1,
    output F2A_B_30_10,
    output F2A_B_30_11,
    output F2A_B_30_12,
    output F2A_B_30_13,
    output F2A_B_30_14,
    output F2A_B_30_15,
    output F2A_B_30_16,
    output F2A_B_30_17,
    output F2A_B_30_2,
    output F2A_B_30_3,
    output F2A_B_30_4,
    output F2A_B_30_5,
    output F2A_B_30_6,
    output F2A_B_30_7,
    output F2A_B_30_8,
    output F2A_B_30_9,
    output F2A_B_31_0,
    output F2A_B_31_1,
    output F2A_B_31_10,
    output F2A_B_31_11,
    output F2A_B_31_2,
    output F2A_B_31_3,
    output F2A_B_31_4,
    output F2A_B_31_5,
    output F2A_B_31_6,
    output F2A_B_31_7,
    output F2A_B_31_8,
    output F2A_B_31_9,
    output F2A_B_32_0,
    output F2A_B_32_1,
    output F2A_B_32_10,
    output F2A_B_32_11,
    output F2A_B_32_12,
    output F2A_B_32_13,
    output F2A_B_32_14,
    output F2A_B_32_15,
    output F2A_B_32_16,
    output F2A_B_32_17,
    output F2A_B_32_2,
    output F2A_B_32_3,
    output F2A_B_32_4,
    output F2A_B_32_5,
    output F2A_B_32_6,
    output F2A_B_32_7,
    output F2A_B_32_8,
    output F2A_B_32_9,
    output F2A_B_3_0,
    output F2A_B_3_1,
    output F2A_B_3_10,
    output F2A_B_3_11,
    output F2A_B_3_2,
    output F2A_B_3_3,
    output F2A_B_3_4,
    output F2A_B_3_5,
    output F2A_B_3_6,
    output F2A_B_3_7,
    output F2A_B_3_8,
    output F2A_B_3_9,
    output F2A_B_4_0,
    output F2A_B_4_1,
    output F2A_B_4_10,
    output F2A_B_4_11,
    output F2A_B_4_12,
    output F2A_B_4_13,
    output F2A_B_4_14,
    output F2A_B_4_15,
    output F2A_B_4_16,
    output F2A_B_4_17,
    output F2A_B_4_2,
    output F2A_B_4_3,
    output F2A_B_4_4,
    output F2A_B_4_5,
    output F2A_B_4_6,
    output F2A_B_4_7,
    output F2A_B_4_8,
    output F2A_B_4_9,
    output F2A_B_5_0,
    output F2A_B_5_1,
    output F2A_B_5_10,
    output F2A_B_5_11,
    output F2A_B_5_2,
    output F2A_B_5_3,
    output F2A_B_5_4,
    output F2A_B_5_5,
    output F2A_B_5_6,
    output F2A_B_5_7,
    output F2A_B_5_8,
    output F2A_B_5_9,
    output F2A_B_6_0,
    output F2A_B_6_1,
    output F2A_B_6_10,
    output F2A_B_6_11,
    output F2A_B_6_12,
    output F2A_B_6_13,
    output F2A_B_6_14,
    output F2A_B_6_15,
    output F2A_B_6_16,
    output F2A_B_6_17,
    output F2A_B_6_2,
    output F2A_B_6_3,
    output F2A_B_6_4,
    output F2A_B_6_5,
    output F2A_B_6_6,
    output F2A_B_6_7,
    output F2A_B_6_8,
    output F2A_B_6_9,
    output F2A_B_7_0,
    output F2A_B_7_1,
    output F2A_B_7_10,
    output F2A_B_7_11,
    output F2A_B_7_2,
    output F2A_B_7_3,
    output F2A_B_7_4,
    output F2A_B_7_5,
    output F2A_B_7_6,
    output F2A_B_7_7,
    output F2A_B_7_8,
    output F2A_B_7_9,
    output F2A_B_8_0,
    output F2A_B_8_1,
    output F2A_B_8_10,
    output F2A_B_8_11,
    output F2A_B_8_12,
    output F2A_B_8_13,
    output F2A_B_8_14,
    output F2A_B_8_15,
    output F2A_B_8_16,
    output F2A_B_8_17,
    output F2A_B_8_2,
    output F2A_B_8_3,
    output F2A_B_8_4,
    output F2A_B_8_5,
    output F2A_B_8_6,
    output F2A_B_8_7,
    output F2A_B_8_8,
    output F2A_B_8_9,
    output F2A_B_9_0,
    output F2A_B_9_1,
    output F2A_B_9_10,
    output F2A_B_9_11,
    output F2A_B_9_2,
    output F2A_B_9_3,
    output F2A_B_9_4,
    output F2A_B_9_5,
    output F2A_B_9_6,
    output F2A_B_9_7,
    output F2A_B_9_8,
    output F2A_B_9_9,
    output F2A_L_10_0,
    output F2A_L_10_1,
    output F2A_L_10_10,
    output F2A_L_10_11,
    output F2A_L_10_12,
    output F2A_L_10_13,
    output F2A_L_10_14,
    output F2A_L_10_15,
    output F2A_L_10_16,
    output F2A_L_10_17,
    output F2A_L_10_2,
    output F2A_L_10_3,
    output F2A_L_10_4,
    output F2A_L_10_5,
    output F2A_L_10_6,
    output F2A_L_10_7,
    output F2A_L_10_8,
    output F2A_L_10_9,
    output F2A_L_11_0,
    output F2A_L_11_1,
    output F2A_L_11_10,
    output F2A_L_11_11,
    output F2A_L_11_2,
    output F2A_L_11_3,
    output F2A_L_11_4,
    output F2A_L_11_5,
    output F2A_L_11_6,
    output F2A_L_11_7,
    output F2A_L_11_8,
    output F2A_L_11_9,
    output F2A_L_12_0,
    output F2A_L_12_1,
    output F2A_L_12_10,
    output F2A_L_12_11,
    output F2A_L_12_12,
    output F2A_L_12_13,
    output F2A_L_12_14,
    output F2A_L_12_15,
    output F2A_L_12_16,
    output F2A_L_12_17,
    output F2A_L_12_2,
    output F2A_L_12_3,
    output F2A_L_12_4,
    output F2A_L_12_5,
    output F2A_L_12_6,
    output F2A_L_12_7,
    output F2A_L_12_8,
    output F2A_L_12_9,
    output F2A_L_13_0,
    output F2A_L_13_1,
    output F2A_L_13_10,
    output F2A_L_13_11,
    output F2A_L_13_2,
    output F2A_L_13_3,
    output F2A_L_13_4,
    output F2A_L_13_5,
    output F2A_L_13_6,
    output F2A_L_13_7,
    output F2A_L_13_8,
    output F2A_L_13_9,
    output F2A_L_14_0,
    output F2A_L_14_1,
    output F2A_L_14_10,
    output F2A_L_14_11,
    output F2A_L_14_12,
    output F2A_L_14_13,
    output F2A_L_14_14,
    output F2A_L_14_15,
    output F2A_L_14_16,
    output F2A_L_14_17,
    output F2A_L_14_2,
    output F2A_L_14_3,
    output F2A_L_14_4,
    output F2A_L_14_5,
    output F2A_L_14_6,
    output F2A_L_14_7,
    output F2A_L_14_8,
    output F2A_L_14_9,
    output F2A_L_15_0,
    output F2A_L_15_1,
    output F2A_L_15_10,
    output F2A_L_15_11,
    output F2A_L_15_2,
    output F2A_L_15_3,
    output F2A_L_15_4,
    output F2A_L_15_5,
    output F2A_L_15_6,
    output F2A_L_15_7,
    output F2A_L_15_8,
    output F2A_L_15_9,
    output F2A_L_16_0,
    output F2A_L_16_1,
    output F2A_L_16_10,
    output F2A_L_16_11,
    output F2A_L_16_12,
    output F2A_L_16_13,
    output F2A_L_16_14,
    output F2A_L_16_15,
    output F2A_L_16_16,
    output F2A_L_16_17,
    output F2A_L_16_2,
    output F2A_L_16_3,
    output F2A_L_16_4,
    output F2A_L_16_5,
    output F2A_L_16_6,
    output F2A_L_16_7,
    output F2A_L_16_8,
    output F2A_L_16_9,
    output F2A_L_17_0,
    output F2A_L_17_1,
    output F2A_L_17_10,
    output F2A_L_17_11,
    output F2A_L_17_2,
    output F2A_L_17_3,
    output F2A_L_17_4,
    output F2A_L_17_5,
    output F2A_L_17_6,
    output F2A_L_17_7,
    output F2A_L_17_8,
    output F2A_L_17_9,
    output F2A_L_18_0,
    output F2A_L_18_1,
    output F2A_L_18_10,
    output F2A_L_18_11,
    output F2A_L_18_12,
    output F2A_L_18_13,
    output F2A_L_18_14,
    output F2A_L_18_15,
    output F2A_L_18_16,
    output F2A_L_18_17,
    output F2A_L_18_2,
    output F2A_L_18_3,
    output F2A_L_18_4,
    output F2A_L_18_5,
    output F2A_L_18_6,
    output F2A_L_18_7,
    output F2A_L_18_8,
    output F2A_L_18_9,
    output F2A_L_19_0,
    output F2A_L_19_1,
    output F2A_L_19_10,
    output F2A_L_19_11,
    output F2A_L_19_2,
    output F2A_L_19_3,
    output F2A_L_19_4,
    output F2A_L_19_5,
    output F2A_L_19_6,
    output F2A_L_19_7,
    output F2A_L_19_8,
    output F2A_L_19_9,
    output F2A_L_1_0,
    output F2A_L_1_1,
    output F2A_L_1_10,
    output F2A_L_1_11,
    output F2A_L_1_2,
    output F2A_L_1_3,
    output F2A_L_1_4,
    output F2A_L_1_5,
    output F2A_L_1_6,
    output F2A_L_1_7,
    output F2A_L_1_8,
    output F2A_L_1_9,
    output F2A_L_20_0,
    output F2A_L_20_1,
    output F2A_L_20_10,
    output F2A_L_20_11,
    output F2A_L_20_12,
    output F2A_L_20_13,
    output F2A_L_20_14,
    output F2A_L_20_15,
    output F2A_L_20_16,
    output F2A_L_20_17,
    output F2A_L_20_2,
    output F2A_L_20_3,
    output F2A_L_20_4,
    output F2A_L_20_5,
    output F2A_L_20_6,
    output F2A_L_20_7,
    output F2A_L_20_8,
    output F2A_L_20_9,
    output F2A_L_21_0,
    output F2A_L_21_1,
    output F2A_L_21_10,
    output F2A_L_21_11,
    output F2A_L_21_2,
    output F2A_L_21_3,
    output F2A_L_21_4,
    output F2A_L_21_5,
    output F2A_L_21_6,
    output F2A_L_21_7,
    output F2A_L_21_8,
    output F2A_L_21_9,
    output F2A_L_22_0,
    output F2A_L_22_1,
    output F2A_L_22_10,
    output F2A_L_22_11,
    output F2A_L_22_12,
    output F2A_L_22_13,
    output F2A_L_22_14,
    output F2A_L_22_15,
    output F2A_L_22_16,
    output F2A_L_22_17,
    output F2A_L_22_2,
    output F2A_L_22_3,
    output F2A_L_22_4,
    output F2A_L_22_5,
    output F2A_L_22_6,
    output F2A_L_22_7,
    output F2A_L_22_8,
    output F2A_L_22_9,
    output F2A_L_23_0,
    output F2A_L_23_1,
    output F2A_L_23_10,
    output F2A_L_23_11,
    output F2A_L_23_2,
    output F2A_L_23_3,
    output F2A_L_23_4,
    output F2A_L_23_5,
    output F2A_L_23_6,
    output F2A_L_23_7,
    output F2A_L_23_8,
    output F2A_L_23_9,
    output F2A_L_24_0,
    output F2A_L_24_1,
    output F2A_L_24_10,
    output F2A_L_24_11,
    output F2A_L_24_12,
    output F2A_L_24_13,
    output F2A_L_24_14,
    output F2A_L_24_15,
    output F2A_L_24_16,
    output F2A_L_24_17,
    output F2A_L_24_2,
    output F2A_L_24_3,
    output F2A_L_24_4,
    output F2A_L_24_5,
    output F2A_L_24_6,
    output F2A_L_24_7,
    output F2A_L_24_8,
    output F2A_L_24_9,
    output F2A_L_25_0,
    output F2A_L_25_1,
    output F2A_L_25_10,
    output F2A_L_25_11,
    output F2A_L_25_2,
    output F2A_L_25_3,
    output F2A_L_25_4,
    output F2A_L_25_5,
    output F2A_L_25_6,
    output F2A_L_25_7,
    output F2A_L_25_8,
    output F2A_L_25_9,
    output F2A_L_26_0,
    output F2A_L_26_1,
    output F2A_L_26_10,
    output F2A_L_26_11,
    output F2A_L_26_12,
    output F2A_L_26_13,
    output F2A_L_26_14,
    output F2A_L_26_15,
    output F2A_L_26_16,
    output F2A_L_26_17,
    output F2A_L_26_2,
    output F2A_L_26_3,
    output F2A_L_26_4,
    output F2A_L_26_5,
    output F2A_L_26_6,
    output F2A_L_26_7,
    output F2A_L_26_8,
    output F2A_L_26_9,
    output F2A_L_27_0,
    output F2A_L_27_1,
    output F2A_L_27_10,
    output F2A_L_27_11,
    output F2A_L_27_2,
    output F2A_L_27_3,
    output F2A_L_27_4,
    output F2A_L_27_5,
    output F2A_L_27_6,
    output F2A_L_27_7,
    output F2A_L_27_8,
    output F2A_L_27_9,
    output F2A_L_28_0,
    output F2A_L_28_1,
    output F2A_L_28_10,
    output F2A_L_28_11,
    output F2A_L_28_12,
    output F2A_L_28_13,
    output F2A_L_28_14,
    output F2A_L_28_15,
    output F2A_L_28_16,
    output F2A_L_28_17,
    output F2A_L_28_2,
    output F2A_L_28_3,
    output F2A_L_28_4,
    output F2A_L_28_5,
    output F2A_L_28_6,
    output F2A_L_28_7,
    output F2A_L_28_8,
    output F2A_L_28_9,
    output F2A_L_29_0,
    output F2A_L_29_1,
    output F2A_L_29_10,
    output F2A_L_29_11,
    output F2A_L_29_2,
    output F2A_L_29_3,
    output F2A_L_29_4,
    output F2A_L_29_5,
    output F2A_L_29_6,
    output F2A_L_29_7,
    output F2A_L_29_8,
    output F2A_L_29_9,
    output F2A_L_2_0,
    output F2A_L_2_1,
    output F2A_L_2_10,
    output F2A_L_2_11,
    output F2A_L_2_12,
    output F2A_L_2_13,
    output F2A_L_2_14,
    output F2A_L_2_15,
    output F2A_L_2_16,
    output F2A_L_2_17,
    output F2A_L_2_2,
    output F2A_L_2_3,
    output F2A_L_2_4,
    output F2A_L_2_5,
    output F2A_L_2_6,
    output F2A_L_2_7,
    output F2A_L_2_8,
    output F2A_L_2_9,
    output F2A_L_30_0,
    output F2A_L_30_1,
    output F2A_L_30_10,
    output F2A_L_30_11,
    output F2A_L_30_12,
    output F2A_L_30_13,
    output F2A_L_30_14,
    output F2A_L_30_15,
    output F2A_L_30_16,
    output F2A_L_30_17,
    output F2A_L_30_2,
    output F2A_L_30_3,
    output F2A_L_30_4,
    output F2A_L_30_5,
    output F2A_L_30_6,
    output F2A_L_30_7,
    output F2A_L_30_8,
    output F2A_L_30_9,
    output F2A_L_31_0,
    output F2A_L_31_1,
    output F2A_L_31_10,
    output F2A_L_31_11,
    output F2A_L_31_2,
    output F2A_L_31_3,
    output F2A_L_31_4,
    output F2A_L_31_5,
    output F2A_L_31_6,
    output F2A_L_31_7,
    output F2A_L_31_8,
    output F2A_L_31_9,
    output F2A_L_32_0,
    output F2A_L_32_1,
    output F2A_L_32_10,
    output F2A_L_32_11,
    output F2A_L_32_12,
    output F2A_L_32_13,
    output F2A_L_32_14,
    output F2A_L_32_15,
    output F2A_L_32_16,
    output F2A_L_32_17,
    output F2A_L_32_2,
    output F2A_L_32_3,
    output F2A_L_32_4,
    output F2A_L_32_5,
    output F2A_L_32_6,
    output F2A_L_32_7,
    output F2A_L_32_8,
    output F2A_L_32_9,
    output F2A_L_3_0,
    output F2A_L_3_1,
    output F2A_L_3_10,
    output F2A_L_3_11,
    output F2A_L_3_2,
    output F2A_L_3_3,
    output F2A_L_3_4,
    output F2A_L_3_5,
    output F2A_L_3_6,
    output F2A_L_3_7,
    output F2A_L_3_8,
    output F2A_L_3_9,
    output F2A_L_4_0,
    output F2A_L_4_1,
    output F2A_L_4_10,
    output F2A_L_4_11,
    output F2A_L_4_12,
    output F2A_L_4_13,
    output F2A_L_4_14,
    output F2A_L_4_15,
    output F2A_L_4_16,
    output F2A_L_4_17,
    output F2A_L_4_2,
    output F2A_L_4_3,
    output F2A_L_4_4,
    output F2A_L_4_5,
    output F2A_L_4_6,
    output F2A_L_4_7,
    output F2A_L_4_8,
    output F2A_L_4_9,
    output F2A_L_5_0,
    output F2A_L_5_1,
    output F2A_L_5_10,
    output F2A_L_5_11,
    output F2A_L_5_2,
    output F2A_L_5_3,
    output F2A_L_5_4,
    output F2A_L_5_5,
    output F2A_L_5_6,
    output F2A_L_5_7,
    output F2A_L_5_8,
    output F2A_L_5_9,
    output F2A_L_6_0,
    output F2A_L_6_1,
    output F2A_L_6_10,
    output F2A_L_6_11,
    output F2A_L_6_12,
    output F2A_L_6_13,
    output F2A_L_6_14,
    output F2A_L_6_15,
    output F2A_L_6_16,
    output F2A_L_6_17,
    output F2A_L_6_2,
    output F2A_L_6_3,
    output F2A_L_6_4,
    output F2A_L_6_5,
    output F2A_L_6_6,
    output F2A_L_6_7,
    output F2A_L_6_8,
    output F2A_L_6_9,
    output F2A_L_7_0,
    output F2A_L_7_1,
    output F2A_L_7_10,
    output F2A_L_7_11,
    output F2A_L_7_2,
    output F2A_L_7_3,
    output F2A_L_7_4,
    output F2A_L_7_5,
    output F2A_L_7_6,
    output F2A_L_7_7,
    output F2A_L_7_8,
    output F2A_L_7_9,
    output F2A_L_8_0,
    output F2A_L_8_1,
    output F2A_L_8_10,
    output F2A_L_8_11,
    output F2A_L_8_12,
    output F2A_L_8_13,
    output F2A_L_8_14,
    output F2A_L_8_15,
    output F2A_L_8_16,
    output F2A_L_8_17,
    output F2A_L_8_2,
    output F2A_L_8_3,
    output F2A_L_8_4,
    output F2A_L_8_5,
    output F2A_L_8_6,
    output F2A_L_8_7,
    output F2A_L_8_8,
    output F2A_L_8_9,
    output F2A_L_9_0,
    output F2A_L_9_1,
    output F2A_L_9_10,
    output F2A_L_9_11,
    output F2A_L_9_2,
    output F2A_L_9_3,
    output F2A_L_9_4,
    output F2A_L_9_5,
    output F2A_L_9_6,
    output F2A_L_9_7,
    output F2A_L_9_8,
    output F2A_L_9_9,
    output F2A_R_10_0,
    output F2A_R_10_1,
    output F2A_R_10_10,
    output F2A_R_10_11,
    output F2A_R_10_12,
    output F2A_R_10_13,
    output F2A_R_10_14,
    output F2A_R_10_15,
    output F2A_R_10_16,
    output F2A_R_10_17,
    output F2A_R_10_2,
    output F2A_R_10_3,
    output F2A_R_10_4,
    output F2A_R_10_5,
    output F2A_R_10_6,
    output F2A_R_10_7,
    output F2A_R_10_8,
    output F2A_R_10_9,
    output F2A_R_11_0,
    output F2A_R_11_1,
    output F2A_R_11_10,
    output F2A_R_11_11,
    output F2A_R_11_2,
    output F2A_R_11_3,
    output F2A_R_11_4,
    output F2A_R_11_5,
    output F2A_R_11_6,
    output F2A_R_11_7,
    output F2A_R_11_8,
    output F2A_R_11_9,
    output F2A_R_12_0,
    output F2A_R_12_1,
    output F2A_R_12_10,
    output F2A_R_12_11,
    output F2A_R_12_12,
    output F2A_R_12_13,
    output F2A_R_12_14,
    output F2A_R_12_15,
    output F2A_R_12_16,
    output F2A_R_12_17,
    output F2A_R_12_2,
    output F2A_R_12_3,
    output F2A_R_12_4,
    output F2A_R_12_5,
    output F2A_R_12_6,
    output F2A_R_12_7,
    output F2A_R_12_8,
    output F2A_R_12_9,
    output F2A_R_13_0,
    output F2A_R_13_1,
    output F2A_R_13_10,
    output F2A_R_13_11,
    output F2A_R_13_2,
    output F2A_R_13_3,
    output F2A_R_13_4,
    output F2A_R_13_5,
    output F2A_R_13_6,
    output F2A_R_13_7,
    output F2A_R_13_8,
    output F2A_R_13_9,
    output F2A_R_14_0,
    output F2A_R_14_1,
    output F2A_R_14_10,
    output F2A_R_14_11,
    output F2A_R_14_12,
    output F2A_R_14_13,
    output F2A_R_14_14,
    output F2A_R_14_15,
    output F2A_R_14_16,
    output F2A_R_14_17,
    output F2A_R_14_2,
    output F2A_R_14_3,
    output F2A_R_14_4,
    output F2A_R_14_5,
    output F2A_R_14_6,
    output F2A_R_14_7,
    output F2A_R_14_8,
    output F2A_R_14_9,
    output F2A_R_15_0,
    output F2A_R_15_1,
    output F2A_R_15_10,
    output F2A_R_15_11,
    output F2A_R_15_2,
    output F2A_R_15_3,
    output F2A_R_15_4,
    output F2A_R_15_5,
    output F2A_R_15_6,
    output F2A_R_15_7,
    output F2A_R_15_8,
    output F2A_R_15_9,
    output F2A_R_16_0,
    output F2A_R_16_1,
    output F2A_R_16_10,
    output F2A_R_16_11,
    output F2A_R_16_12,
    output F2A_R_16_13,
    output F2A_R_16_14,
    output F2A_R_16_15,
    output F2A_R_16_16,
    output F2A_R_16_17,
    output F2A_R_16_2,
    output F2A_R_16_3,
    output F2A_R_16_4,
    output F2A_R_16_5,
    output F2A_R_16_6,
    output F2A_R_16_7,
    output F2A_R_16_8,
    output F2A_R_16_9,
    output F2A_R_17_0,
    output F2A_R_17_1,
    output F2A_R_17_10,
    output F2A_R_17_11,
    output F2A_R_17_2,
    output F2A_R_17_3,
    output F2A_R_17_4,
    output F2A_R_17_5,
    output F2A_R_17_6,
    output F2A_R_17_7,
    output F2A_R_17_8,
    output F2A_R_17_9,
    output F2A_R_18_0,
    output F2A_R_18_1,
    output F2A_R_18_10,
    output F2A_R_18_11,
    output F2A_R_18_12,
    output F2A_R_18_13,
    output F2A_R_18_14,
    output F2A_R_18_15,
    output F2A_R_18_16,
    output F2A_R_18_17,
    output F2A_R_18_2,
    output F2A_R_18_3,
    output F2A_R_18_4,
    output F2A_R_18_5,
    output F2A_R_18_6,
    output F2A_R_18_7,
    output F2A_R_18_8,
    output F2A_R_18_9,
    output F2A_R_19_0,
    output F2A_R_19_1,
    output F2A_R_19_10,
    output F2A_R_19_11,
    output F2A_R_19_2,
    output F2A_R_19_3,
    output F2A_R_19_4,
    output F2A_R_19_5,
    output F2A_R_19_6,
    output F2A_R_19_7,
    output F2A_R_19_8,
    output F2A_R_19_9,
    output F2A_R_1_0,
    output F2A_R_1_1,
    output F2A_R_1_10,
    output F2A_R_1_11,
    output F2A_R_1_2,
    output F2A_R_1_3,
    output F2A_R_1_4,
    output F2A_R_1_5,
    output F2A_R_1_6,
    output F2A_R_1_7,
    output F2A_R_1_8,
    output F2A_R_1_9,
    output F2A_R_20_0,
    output F2A_R_20_1,
    output F2A_R_20_10,
    output F2A_R_20_11,
    output F2A_R_20_12,
    output F2A_R_20_13,
    output F2A_R_20_14,
    output F2A_R_20_15,
    output F2A_R_20_16,
    output F2A_R_20_17,
    output F2A_R_20_2,
    output F2A_R_20_3,
    output F2A_R_20_4,
    output F2A_R_20_5,
    output F2A_R_20_6,
    output F2A_R_20_7,
    output F2A_R_20_8,
    output F2A_R_20_9,
    output F2A_R_21_0,
    output F2A_R_21_1,
    output F2A_R_21_10,
    output F2A_R_21_11,
    output F2A_R_21_2,
    output F2A_R_21_3,
    output F2A_R_21_4,
    output F2A_R_21_5,
    output F2A_R_21_6,
    output F2A_R_21_7,
    output F2A_R_21_8,
    output F2A_R_21_9,
    output F2A_R_22_0,
    output F2A_R_22_1,
    output F2A_R_22_10,
    output F2A_R_22_11,
    output F2A_R_22_12,
    output F2A_R_22_13,
    output F2A_R_22_14,
    output F2A_R_22_15,
    output F2A_R_22_16,
    output F2A_R_22_17,
    output F2A_R_22_2,
    output F2A_R_22_3,
    output F2A_R_22_4,
    output F2A_R_22_5,
    output F2A_R_22_6,
    output F2A_R_22_7,
    output F2A_R_22_8,
    output F2A_R_22_9,
    output F2A_R_23_0,
    output F2A_R_23_1,
    output F2A_R_23_10,
    output F2A_R_23_11,
    output F2A_R_23_2,
    output F2A_R_23_3,
    output F2A_R_23_4,
    output F2A_R_23_5,
    output F2A_R_23_6,
    output F2A_R_23_7,
    output F2A_R_23_8,
    output F2A_R_23_9,
    output F2A_R_24_0,
    output F2A_R_24_1,
    output F2A_R_24_10,
    output F2A_R_24_11,
    output F2A_R_24_12,
    output F2A_R_24_13,
    output F2A_R_24_14,
    output F2A_R_24_15,
    output F2A_R_24_16,
    output F2A_R_24_17,
    output F2A_R_24_2,
    output F2A_R_24_3,
    output F2A_R_24_4,
    output F2A_R_24_5,
    output F2A_R_24_6,
    output F2A_R_24_7,
    output F2A_R_24_8,
    output F2A_R_24_9,
    output F2A_R_25_0,
    output F2A_R_25_1,
    output F2A_R_25_10,
    output F2A_R_25_11,
    output F2A_R_25_2,
    output F2A_R_25_3,
    output F2A_R_25_4,
    output F2A_R_25_5,
    output F2A_R_25_6,
    output F2A_R_25_7,
    output F2A_R_25_8,
    output F2A_R_25_9,
    output F2A_R_26_0,
    output F2A_R_26_1,
    output F2A_R_26_10,
    output F2A_R_26_11,
    output F2A_R_26_12,
    output F2A_R_26_13,
    output F2A_R_26_14,
    output F2A_R_26_15,
    output F2A_R_26_16,
    output F2A_R_26_17,
    output F2A_R_26_2,
    output F2A_R_26_3,
    output F2A_R_26_4,
    output F2A_R_26_5,
    output F2A_R_26_6,
    output F2A_R_26_7,
    output F2A_R_26_8,
    output F2A_R_26_9,
    output F2A_R_27_0,
    output F2A_R_27_1,
    output F2A_R_27_10,
    output F2A_R_27_11,
    output F2A_R_27_2,
    output F2A_R_27_3,
    output F2A_R_27_4,
    output F2A_R_27_5,
    output F2A_R_27_6,
    output F2A_R_27_7,
    output F2A_R_27_8,
    output F2A_R_27_9,
    output F2A_R_28_0,
    output F2A_R_28_1,
    output F2A_R_28_10,
    output F2A_R_28_11,
    output F2A_R_28_12,
    output F2A_R_28_13,
    output F2A_R_28_14,
    output F2A_R_28_15,
    output F2A_R_28_16,
    output F2A_R_28_17,
    output F2A_R_28_2,
    output F2A_R_28_3,
    output F2A_R_28_4,
    output F2A_R_28_5,
    output F2A_R_28_6,
    output F2A_R_28_7,
    output F2A_R_28_8,
    output F2A_R_28_9,
    output F2A_R_29_0,
    output F2A_R_29_1,
    output F2A_R_29_10,
    output F2A_R_29_11,
    output F2A_R_29_2,
    output F2A_R_29_3,
    output F2A_R_29_4,
    output F2A_R_29_5,
    output F2A_R_29_6,
    output F2A_R_29_7,
    output F2A_R_29_8,
    output F2A_R_29_9,
    output F2A_R_2_0,
    output F2A_R_2_1,
    output F2A_R_2_10,
    output F2A_R_2_11,
    output F2A_R_2_12,
    output F2A_R_2_13,
    output F2A_R_2_14,
    output F2A_R_2_15,
    output F2A_R_2_16,
    output F2A_R_2_17,
    output F2A_R_2_2,
    output F2A_R_2_3,
    output F2A_R_2_4,
    output F2A_R_2_5,
    output F2A_R_2_6,
    output F2A_R_2_7,
    output F2A_R_2_8,
    output F2A_R_2_9,
    output F2A_R_30_0,
    output F2A_R_30_1,
    output F2A_R_30_10,
    output F2A_R_30_11,
    output F2A_R_30_12,
    output F2A_R_30_13,
    output F2A_R_30_14,
    output F2A_R_30_15,
    output F2A_R_30_16,
    output F2A_R_30_17,
    output F2A_R_30_2,
    output F2A_R_30_3,
    output F2A_R_30_4,
    output F2A_R_30_5,
    output F2A_R_30_6,
    output F2A_R_30_7,
    output F2A_R_30_8,
    output F2A_R_30_9,
    output F2A_R_31_0,
    output F2A_R_31_1,
    output F2A_R_31_10,
    output F2A_R_31_11,
    output F2A_R_31_2,
    output F2A_R_31_3,
    output F2A_R_31_4,
    output F2A_R_31_5,
    output F2A_R_31_6,
    output F2A_R_31_7,
    output F2A_R_31_8,
    output F2A_R_31_9,
    output F2A_R_32_0,
    output F2A_R_32_1,
    output F2A_R_32_10,
    output F2A_R_32_11,
    output F2A_R_32_12,
    output F2A_R_32_13,
    output F2A_R_32_14,
    output F2A_R_32_15,
    output F2A_R_32_16,
    output F2A_R_32_17,
    output F2A_R_32_2,
    output F2A_R_32_3,
    output F2A_R_32_4,
    output F2A_R_32_5,
    output F2A_R_32_6,
    output F2A_R_32_7,
    output F2A_R_32_8,
    output F2A_R_32_9,
    output F2A_R_3_0,
    output F2A_R_3_1,
    output F2A_R_3_10,
    output F2A_R_3_11,
    output F2A_R_3_2,
    output F2A_R_3_3,
    output F2A_R_3_4,
    output F2A_R_3_5,
    output F2A_R_3_6,
    output F2A_R_3_7,
    output F2A_R_3_8,
    output F2A_R_3_9,
    output F2A_R_4_0,
    output F2A_R_4_1,
    output F2A_R_4_10,
    output F2A_R_4_11,
    output F2A_R_4_12,
    output F2A_R_4_13,
    output F2A_R_4_14,
    output F2A_R_4_15,
    output F2A_R_4_16,
    output F2A_R_4_17,
    output F2A_R_4_2,
    output F2A_R_4_3,
    output F2A_R_4_4,
    output F2A_R_4_5,
    output F2A_R_4_6,
    output F2A_R_4_7,
    output F2A_R_4_8,
    output F2A_R_4_9,
    output F2A_R_5_0,
    output F2A_R_5_1,
    output F2A_R_5_10,
    output F2A_R_5_11,
    output F2A_R_5_2,
    output F2A_R_5_3,
    output F2A_R_5_4,
    output F2A_R_5_5,
    output F2A_R_5_6,
    output F2A_R_5_7,
    output F2A_R_5_8,
    output F2A_R_5_9,
    output F2A_R_6_0,
    output F2A_R_6_1,
    output F2A_R_6_10,
    output F2A_R_6_11,
    output F2A_R_6_12,
    output F2A_R_6_13,
    output F2A_R_6_14,
    output F2A_R_6_15,
    output F2A_R_6_16,
    output F2A_R_6_17,
    output F2A_R_6_2,
    output F2A_R_6_3,
    output F2A_R_6_4,
    output F2A_R_6_5,
    output F2A_R_6_6,
    output F2A_R_6_7,
    output F2A_R_6_8,
    output F2A_R_6_9,
    output F2A_R_7_0,
    output F2A_R_7_1,
    output F2A_R_7_10,
    output F2A_R_7_11,
    output F2A_R_7_2,
    output F2A_R_7_3,
    output F2A_R_7_4,
    output F2A_R_7_5,
    output F2A_R_7_6,
    output F2A_R_7_7,
    output F2A_R_7_8,
    output F2A_R_7_9,
    output F2A_R_8_0,
    output F2A_R_8_1,
    output F2A_R_8_10,
    output F2A_R_8_11,
    output F2A_R_8_12,
    output F2A_R_8_13,
    output F2A_R_8_14,
    output F2A_R_8_15,
    output F2A_R_8_16,
    output F2A_R_8_17,
    output F2A_R_8_2,
    output F2A_R_8_3,
    output F2A_R_8_4,
    output F2A_R_8_5,
    output F2A_R_8_6,
    output F2A_R_8_7,
    output F2A_R_8_8,
    output F2A_R_8_9,
    output F2A_R_9_0,
    output F2A_R_9_1,
    output F2A_R_9_10,
    output F2A_R_9_11,
    output F2A_R_9_2,
    output F2A_R_9_3,
    output F2A_R_9_4,
    output F2A_R_9_5,
    output F2A_R_9_6,
    output F2A_R_9_7,
    output F2A_R_9_8,
    output F2A_R_9_9,
    output F2A_T_10_0,
    output F2A_T_10_1,
    output F2A_T_10_10,
    output F2A_T_10_11,
    output F2A_T_10_12,
    output F2A_T_10_13,
    output F2A_T_10_14,
    output F2A_T_10_15,
    output F2A_T_10_16,
    output F2A_T_10_17,
    output F2A_T_10_2,
    output F2A_T_10_3,
    output F2A_T_10_4,
    output F2A_T_10_5,
    output F2A_T_10_6,
    output F2A_T_10_7,
    output F2A_T_10_8,
    output F2A_T_10_9,
    output F2A_T_11_0,
    output F2A_T_11_1,
    output F2A_T_11_10,
    output F2A_T_11_11,
    output F2A_T_11_2,
    output F2A_T_11_3,
    output F2A_T_11_4,
    output F2A_T_11_5,
    output F2A_T_11_6,
    output F2A_T_11_7,
    output F2A_T_11_8,
    output F2A_T_11_9,
    output F2A_T_12_0,
    output F2A_T_12_1,
    output F2A_T_12_10,
    output F2A_T_12_11,
    output F2A_T_12_12,
    output F2A_T_12_13,
    output F2A_T_12_14,
    output F2A_T_12_15,
    output F2A_T_12_16,
    output F2A_T_12_17,
    output F2A_T_12_2,
    output F2A_T_12_3,
    output F2A_T_12_4,
    output F2A_T_12_5,
    output F2A_T_12_6,
    output F2A_T_12_7,
    output F2A_T_12_8,
    output F2A_T_12_9,
    output F2A_T_13_0,
    output F2A_T_13_1,
    output F2A_T_13_10,
    output F2A_T_13_11,
    output F2A_T_13_2,
    output F2A_T_13_3,
    output F2A_T_13_4,
    output F2A_T_13_5,
    output F2A_T_13_6,
    output F2A_T_13_7,
    output F2A_T_13_8,
    output F2A_T_13_9,
    output F2A_T_14_0,
    output F2A_T_14_1,
    output F2A_T_14_10,
    output F2A_T_14_11,
    output F2A_T_14_12,
    output F2A_T_14_13,
    output F2A_T_14_14,
    output F2A_T_14_15,
    output F2A_T_14_16,
    output F2A_T_14_17,
    output F2A_T_14_2,
    output F2A_T_14_3,
    output F2A_T_14_4,
    output F2A_T_14_5,
    output F2A_T_14_6,
    output F2A_T_14_7,
    output F2A_T_14_8,
    output F2A_T_14_9,
    output F2A_T_15_0,
    output F2A_T_15_1,
    output F2A_T_15_10,
    output F2A_T_15_11,
    output F2A_T_15_2,
    output F2A_T_15_3,
    output F2A_T_15_4,
    output F2A_T_15_5,
    output F2A_T_15_6,
    output F2A_T_15_7,
    output F2A_T_15_8,
    output F2A_T_15_9,
    output F2A_T_16_0,
    output F2A_T_16_1,
    output F2A_T_16_10,
    output F2A_T_16_11,
    output F2A_T_16_12,
    output F2A_T_16_13,
    output F2A_T_16_17,
    output F2A_T_16_2,
    output F2A_T_16_3,
    output F2A_T_16_4,
    output F2A_T_16_5,
    output F2A_T_16_6,
    output F2A_T_16_7,
    output F2A_T_16_8,
    output F2A_T_16_9,
    output F2A_T_17_0,
    output F2A_T_17_1,
    output F2A_T_17_10,
    output F2A_T_17_11,
    output F2A_T_17_2,
    output F2A_T_17_3,
    output F2A_T_17_4,
    output F2A_T_17_5,
    output F2A_T_17_6,
    output F2A_T_17_7,
    output F2A_T_17_8,
    output F2A_T_17_9,
    output F2A_T_18_0,
    output F2A_T_18_1,
    output F2A_T_18_10,
    output F2A_T_18_11,
    output F2A_T_18_12,
    output F2A_T_18_13,
    output F2A_T_18_14,
    output F2A_T_18_15,
    output F2A_T_18_16,
    output F2A_T_18_17,
    output F2A_T_18_2,
    output F2A_T_18_3,
    output F2A_T_18_4,
    output F2A_T_18_5,
    output F2A_T_18_6,
    output F2A_T_18_7,
    output F2A_T_18_8,
    output F2A_T_18_9,
    output F2A_T_19_0,
    output F2A_T_19_1,
    output F2A_T_19_10,
    output F2A_T_19_11,
    output F2A_T_19_2,
    output F2A_T_19_3,
    output F2A_T_19_4,
    output F2A_T_19_5,
    output F2A_T_19_6,
    output F2A_T_19_7,
    output F2A_T_19_8,
    output F2A_T_19_9,
    output F2A_T_1_0,
    output F2A_T_1_1,
    output F2A_T_1_10,
    output F2A_T_1_11,
    output F2A_T_1_2,
    output F2A_T_1_3,
    output F2A_T_1_4,
    output F2A_T_1_5,
    output F2A_T_1_6,
    output F2A_T_1_7,
    output F2A_T_1_8,
    output F2A_T_1_9,
    output F2A_T_20_0,
    output F2A_T_20_1,
    output F2A_T_20_10,
    output F2A_T_20_11,
    output F2A_T_20_12,
    output F2A_T_20_13,
    output F2A_T_20_14,
    output F2A_T_20_15,
    output F2A_T_20_16,
    output F2A_T_20_17,
    output F2A_T_20_2,
    output F2A_T_20_3,
    output F2A_T_20_4,
    output F2A_T_20_5,
    output F2A_T_20_6,
    output F2A_T_20_7,
    output F2A_T_20_8,
    output F2A_T_20_9,
    output F2A_T_21_0,
    output F2A_T_21_1,
    output F2A_T_21_10,
    output F2A_T_21_11,
    output F2A_T_21_2,
    output F2A_T_21_3,
    output F2A_T_21_4,
    output F2A_T_21_5,
    output F2A_T_21_6,
    output F2A_T_21_7,
    output F2A_T_21_8,
    output F2A_T_21_9,
    output F2A_T_22_0,
    output F2A_T_22_1,
    output F2A_T_22_10,
    output F2A_T_22_11,
    output F2A_T_22_12,
    output F2A_T_22_13,
    output F2A_T_22_14,
    output F2A_T_22_15,
    output F2A_T_22_16,
    output F2A_T_22_17,
    output F2A_T_22_2,
    output F2A_T_22_3,
    output F2A_T_22_4,
    output F2A_T_22_5,
    output F2A_T_22_6,
    output F2A_T_22_7,
    output F2A_T_22_8,
    output F2A_T_22_9,
    output F2A_T_23_0,
    output F2A_T_23_1,
    output F2A_T_23_10,
    output F2A_T_23_11,
    output F2A_T_23_2,
    output F2A_T_23_3,
    output F2A_T_23_4,
    output F2A_T_23_5,
    output F2A_T_23_6,
    output F2A_T_23_7,
    output F2A_T_23_8,
    output F2A_T_23_9,
    output F2A_T_24_0,
    output F2A_T_24_1,
    output F2A_T_24_10,
    output F2A_T_24_11,
    output F2A_T_24_12,
    output F2A_T_24_13,
    output F2A_T_24_14,
    output F2A_T_24_15,
    output F2A_T_24_16,
    output F2A_T_24_17,
    output F2A_T_24_2,
    output F2A_T_24_3,
    output F2A_T_24_4,
    output F2A_T_24_5,
    output F2A_T_24_6,
    output F2A_T_24_7,
    output F2A_T_24_8,
    output F2A_T_24_9,
    output F2A_T_25_0,
    output F2A_T_25_1,
    output F2A_T_25_10,
    output F2A_T_25_11,
    output F2A_T_25_2,
    output F2A_T_25_3,
    output F2A_T_25_4,
    output F2A_T_25_5,
    output F2A_T_25_6,
    output F2A_T_25_7,
    output F2A_T_25_8,
    output F2A_T_25_9,
    output F2A_T_26_0,
    output F2A_T_26_1,
    output F2A_T_26_10,
    output F2A_T_26_11,
    output F2A_T_26_12,
    output F2A_T_26_13,
    output F2A_T_26_14,
    output F2A_T_26_15,
    output F2A_T_26_16,
    output F2A_T_26_17,
    output F2A_T_26_2,
    output F2A_T_26_3,
    output F2A_T_26_4,
    output F2A_T_26_5,
    output F2A_T_26_6,
    output F2A_T_26_7,
    output F2A_T_26_8,
    output F2A_T_26_9,
    output F2A_T_27_0,
    output F2A_T_27_1,
    output F2A_T_27_10,
    output F2A_T_27_11,
    output F2A_T_27_2,
    output F2A_T_27_3,
    output F2A_T_27_4,
    output F2A_T_27_5,
    output F2A_T_27_6,
    output F2A_T_27_7,
    output F2A_T_27_8,
    output F2A_T_27_9,
    output F2A_T_28_0,
    output F2A_T_28_1,
    output F2A_T_28_10,
    output F2A_T_28_11,
    output F2A_T_28_12,
    output F2A_T_28_13,
    output F2A_T_28_14,
    output F2A_T_28_15,
    output F2A_T_28_16,
    output F2A_T_28_17,
    output F2A_T_28_2,
    output F2A_T_28_3,
    output F2A_T_28_4,
    output F2A_T_28_5,
    output F2A_T_28_6,
    output F2A_T_28_7,
    output F2A_T_28_8,
    output F2A_T_28_9,
    output F2A_T_29_0,
    output F2A_T_29_1,
    output F2A_T_29_10,
    output F2A_T_29_11,
    output F2A_T_29_2,
    output F2A_T_29_3,
    output F2A_T_29_4,
    output F2A_T_29_5,
    output F2A_T_29_6,
    output F2A_T_29_7,
    output F2A_T_29_8,
    output F2A_T_29_9,
    output F2A_T_2_0,
    output F2A_T_2_1,
    output F2A_T_2_10,
    output F2A_T_2_11,
    output F2A_T_2_12,
    output F2A_T_2_13,
    output F2A_T_2_14,
    output F2A_T_2_15,
    output F2A_T_2_16,
    output F2A_T_2_17,
    output F2A_T_2_2,
    output F2A_T_2_3,
    output F2A_T_2_4,
    output F2A_T_2_5,
    output F2A_T_2_6,
    output F2A_T_2_7,
    output F2A_T_2_8,
    output F2A_T_2_9,
    output F2A_T_30_0,
    output F2A_T_30_1,
    output F2A_T_30_10,
    output F2A_T_30_11,
    output F2A_T_30_12,
    output F2A_T_30_13,
    output F2A_T_30_14,
    output F2A_T_30_15,
    output F2A_T_30_16,
    output F2A_T_30_17,
    output F2A_T_30_2,
    output F2A_T_30_3,
    output F2A_T_30_4,
    output F2A_T_30_5,
    output F2A_T_30_6,
    output F2A_T_30_7,
    output F2A_T_30_8,
    output F2A_T_30_9,
    output F2A_T_31_0,
    output F2A_T_31_1,
    output F2A_T_31_10,
    output F2A_T_31_11,
    output F2A_T_31_2,
    output F2A_T_31_3,
    output F2A_T_31_4,
    output F2A_T_31_5,
    output F2A_T_31_6,
    output F2A_T_31_7,
    output F2A_T_31_8,
    output F2A_T_31_9,
    output F2A_T_32_0,
    output F2A_T_32_1,
    output F2A_T_32_10,
    output F2A_T_32_11,
    output F2A_T_32_12,
    output F2A_T_32_13,
    output F2A_T_32_14,
    output F2A_T_32_15,
    output F2A_T_32_16,
    output F2A_T_32_17,
    output F2A_T_32_2,
    output F2A_T_32_3,
    output F2A_T_32_4,
    output F2A_T_32_5,
    output F2A_T_32_6,
    output F2A_T_32_7,
    output F2A_T_32_8,
    output F2A_T_32_9,
    output F2A_T_3_0,
    output F2A_T_3_1,
    output F2A_T_3_10,
    output F2A_T_3_11,
    output F2A_T_3_2,
    output F2A_T_3_3,
    output F2A_T_3_4,
    output F2A_T_3_5,
    output F2A_T_3_6,
    output F2A_T_3_7,
    output F2A_T_3_8,
    output F2A_T_3_9,
    output F2A_T_4_0,
    output F2A_T_4_1,
    output F2A_T_4_10,
    output F2A_T_4_11,
    output F2A_T_4_12,
    output F2A_T_4_13,
    output F2A_T_4_14,
    output F2A_T_4_15,
    output F2A_T_4_16,
    output F2A_T_4_17,
    output F2A_T_4_2,
    output F2A_T_4_3,
    output F2A_T_4_4,
    output F2A_T_4_5,
    output F2A_T_4_6,
    output F2A_T_4_7,
    output F2A_T_4_8,
    output F2A_T_4_9,
    output F2A_T_5_0,
    output F2A_T_5_1,
    output F2A_T_5_10,
    output F2A_T_5_11,
    output F2A_T_5_2,
    output F2A_T_5_3,
    output F2A_T_5_4,
    output F2A_T_5_5,
    output F2A_T_5_6,
    output F2A_T_5_7,
    output F2A_T_5_8,
    output F2A_T_5_9,
    output F2A_T_6_0,
    output F2A_T_6_1,
    output F2A_T_6_10,
    output F2A_T_6_11,
    output F2A_T_6_12,
    output F2A_T_6_13,
    output F2A_T_6_14,
    output F2A_T_6_15,
    output F2A_T_6_16,
    output F2A_T_6_17,
    output F2A_T_6_2,
    output F2A_T_6_3,
    output F2A_T_6_4,
    output F2A_T_6_5,
    output F2A_T_6_6,
    output F2A_T_6_7,
    output F2A_T_6_8,
    output F2A_T_6_9,
    output F2A_T_7_0,
    output F2A_T_7_1,
    output F2A_T_7_10,
    output F2A_T_7_11,
    output F2A_T_7_2,
    output F2A_T_7_3,
    output F2A_T_7_4,
    output F2A_T_7_5,
    output F2A_T_7_6,
    output F2A_T_7_7,
    output F2A_T_7_8,
    output F2A_T_7_9,
    output F2A_T_8_0,
    output F2A_T_8_1,
    output F2A_T_8_10,
    output F2A_T_8_11,
    output F2A_T_8_12,
    output F2A_T_8_13,
    output F2A_T_8_14,
    output F2A_T_8_15,
    output F2A_T_8_16,
    output F2A_T_8_17,
    output F2A_T_8_2,
    output F2A_T_8_3,
    output F2A_T_8_4,
    output F2A_T_8_5,
    output F2A_T_8_6,
    output F2A_T_8_7,
    output F2A_T_8_8,
    output F2A_T_8_9,
    output F2A_T_9_0,
    output F2A_T_9_1,
    output F2A_T_9_10,
    output F2A_T_9_11,
    output F2A_T_9_2,
    output F2A_T_9_3,
    output F2A_T_9_4,
    output F2A_T_9_5,
    output F2A_T_9_6,
    output F2A_T_9_7,
    output F2A_T_9_8,
    output F2A_T_9_9,
    output F2Adef_B_10_0,
    output F2Adef_B_10_1,
    output F2Adef_B_10_2,
    output F2Adef_B_10_3,
    output F2Adef_B_10_4,
    output F2Adef_B_10_5,
    output F2Adef_B_10_6,
    output F2Adef_B_11_0,
    output F2Adef_B_11_1,
    output F2Adef_B_11_2,
    output F2Adef_B_11_3,
    output F2Adef_B_12_0,
    output F2Adef_B_12_1,
    output F2Adef_B_12_2,
    output F2Adef_B_12_3,
    output F2Adef_B_12_4,
    output F2Adef_B_12_5,
    output F2Adef_B_12_6,
    output F2Adef_B_13_0,
    output F2Adef_B_13_1,
    output F2Adef_B_13_2,
    output F2Adef_B_13_3,
    output F2Adef_B_14_0,
    output F2Adef_B_14_1,
    output F2Adef_B_14_2,
    output F2Adef_B_14_3,
    output F2Adef_B_14_4,
    output F2Adef_B_14_5,
    output F2Adef_B_14_6,
    output F2Adef_B_15_0,
    output F2Adef_B_15_1,
    output F2Adef_B_15_2,
    output F2Adef_B_15_3,
    output F2Adef_B_16_0,
    output F2Adef_B_16_1,
    output F2Adef_B_16_2,
    output F2Adef_B_16_3,
    output F2Adef_B_16_4,
    output F2Adef_B_16_5,
    output F2Adef_B_16_6,
    output F2Adef_B_17_0,
    output F2Adef_B_17_1,
    output F2Adef_B_17_2,
    output F2Adef_B_17_3,
    output F2Adef_B_18_0,
    output F2Adef_B_18_1,
    output F2Adef_B_18_2,
    output F2Adef_B_18_3,
    output F2Adef_B_18_4,
    output F2Adef_B_18_5,
    output F2Adef_B_18_6,
    output F2Adef_B_19_0,
    output F2Adef_B_19_1,
    output F2Adef_B_19_2,
    output F2Adef_B_19_3,
    output F2Adef_B_1_0,
    output F2Adef_B_1_1,
    output F2Adef_B_1_2,
    output F2Adef_B_1_3,
    output F2Adef_B_20_0,
    output F2Adef_B_20_1,
    output F2Adef_B_20_2,
    output F2Adef_B_20_3,
    output F2Adef_B_20_4,
    output F2Adef_B_20_5,
    output F2Adef_B_20_6,
    output F2Adef_B_21_0,
    output F2Adef_B_21_1,
    output F2Adef_B_21_2,
    output F2Adef_B_21_3,
    output F2Adef_B_22_0,
    output F2Adef_B_22_1,
    output F2Adef_B_22_2,
    output F2Adef_B_22_3,
    output F2Adef_B_22_4,
    output F2Adef_B_22_5,
    output F2Adef_B_22_6,
    output F2Adef_B_23_0,
    output F2Adef_B_23_1,
    output F2Adef_B_23_2,
    output F2Adef_B_23_3,
    output F2Adef_B_24_0,
    output F2Adef_B_24_1,
    output F2Adef_B_24_2,
    output F2Adef_B_24_3,
    output F2Adef_B_24_4,
    output F2Adef_B_24_5,
    output F2Adef_B_24_6,
    output F2Adef_B_25_0,
    output F2Adef_B_25_1,
    output F2Adef_B_25_2,
    output F2Adef_B_25_3,
    output F2Adef_B_26_0,
    output F2Adef_B_26_1,
    output F2Adef_B_26_2,
    output F2Adef_B_26_3,
    output F2Adef_B_26_4,
    output F2Adef_B_26_5,
    output F2Adef_B_26_6,
    output F2Adef_B_27_0,
    output F2Adef_B_27_1,
    output F2Adef_B_27_2,
    output F2Adef_B_27_3,
    output F2Adef_B_28_0,
    output F2Adef_B_28_1,
    output F2Adef_B_28_2,
    output F2Adef_B_28_3,
    output F2Adef_B_28_4,
    output F2Adef_B_28_5,
    output F2Adef_B_28_6,
    output F2Adef_B_29_0,
    output F2Adef_B_29_1,
    output F2Adef_B_29_2,
    output F2Adef_B_29_3,
    output F2Adef_B_2_0,
    output F2Adef_B_2_1,
    output F2Adef_B_2_2,
    output F2Adef_B_2_3,
    output F2Adef_B_2_4,
    output F2Adef_B_2_5,
    output F2Adef_B_2_6,
    output F2Adef_B_30_0,
    output F2Adef_B_30_1,
    output F2Adef_B_30_2,
    output F2Adef_B_30_3,
    output F2Adef_B_30_4,
    output F2Adef_B_30_5,
    output F2Adef_B_30_6,
    output F2Adef_B_31_0,
    output F2Adef_B_31_1,
    output F2Adef_B_31_2,
    output F2Adef_B_31_3,
    output F2Adef_B_32_0,
    output F2Adef_B_32_1,
    output F2Adef_B_32_2,
    output F2Adef_B_32_3,
    output F2Adef_B_32_4,
    output F2Adef_B_32_5,
    output F2Adef_B_32_6,
    output F2Adef_B_3_0,
    output F2Adef_B_3_1,
    output F2Adef_B_3_2,
    output F2Adef_B_3_3,
    output F2Adef_B_4_0,
    output F2Adef_B_4_1,
    output F2Adef_B_4_2,
    output F2Adef_B_4_3,
    output F2Adef_B_4_4,
    output F2Adef_B_4_5,
    output F2Adef_B_4_6,
    output F2Adef_B_5_0,
    output F2Adef_B_5_1,
    output F2Adef_B_5_2,
    output F2Adef_B_5_3,
    output F2Adef_B_6_0,
    output F2Adef_B_6_1,
    output F2Adef_B_6_2,
    output F2Adef_B_6_3,
    output F2Adef_B_6_4,
    output F2Adef_B_6_5,
    output F2Adef_B_6_6,
    output F2Adef_B_7_0,
    output F2Adef_B_7_1,
    output F2Adef_B_7_2,
    output F2Adef_B_7_3,
    output F2Adef_B_8_0,
    output F2Adef_B_8_1,
    output F2Adef_B_8_2,
    output F2Adef_B_8_3,
    output F2Adef_B_8_4,
    output F2Adef_B_8_5,
    output F2Adef_B_8_6,
    output F2Adef_B_9_0,
    output F2Adef_B_9_1,
    output F2Adef_B_9_2,
    output F2Adef_B_9_3,
    output F2Adef_L_10_0,
    output F2Adef_L_10_1,
    output F2Adef_L_10_2,
    output F2Adef_L_10_3,
    output F2Adef_L_10_4,
    output F2Adef_L_10_5,
    output F2Adef_L_10_6,
    output F2Adef_L_11_0,
    output F2Adef_L_11_1,
    output F2Adef_L_11_2,
    output F2Adef_L_11_3,
    output F2Adef_L_12_0,
    output F2Adef_L_12_1,
    output F2Adef_L_12_2,
    output F2Adef_L_12_3,
    output F2Adef_L_12_4,
    output F2Adef_L_12_5,
    output F2Adef_L_12_6,
    output F2Adef_L_13_0,
    output F2Adef_L_13_1,
    output F2Adef_L_13_2,
    output F2Adef_L_13_3,
    output F2Adef_L_14_0,
    output F2Adef_L_14_1,
    output F2Adef_L_14_2,
    output F2Adef_L_14_3,
    output F2Adef_L_14_4,
    output F2Adef_L_14_5,
    output F2Adef_L_14_6,
    output F2Adef_L_15_0,
    output F2Adef_L_15_1,
    output F2Adef_L_15_2,
    output F2Adef_L_15_3,
    output F2Adef_L_16_0,
    output F2Adef_L_16_1,
    output F2Adef_L_16_2,
    output F2Adef_L_16_3,
    output F2Adef_L_16_4,
    output F2Adef_L_16_5,
    output F2Adef_L_16_6,
    output F2Adef_L_17_0,
    output F2Adef_L_17_1,
    output F2Adef_L_17_2,
    output F2Adef_L_17_3,
    output F2Adef_L_18_0,
    output F2Adef_L_18_1,
    output F2Adef_L_18_2,
    output F2Adef_L_18_3,
    output F2Adef_L_18_4,
    output F2Adef_L_18_5,
    output F2Adef_L_18_6,
    output F2Adef_L_19_0,
    output F2Adef_L_19_1,
    output F2Adef_L_19_2,
    output F2Adef_L_19_3,
    output F2Adef_L_1_0,
    output F2Adef_L_1_1,
    output F2Adef_L_1_2,
    output F2Adef_L_1_3,
    output F2Adef_L_20_0,
    output F2Adef_L_20_1,
    output F2Adef_L_20_2,
    output F2Adef_L_20_3,
    output F2Adef_L_20_4,
    output F2Adef_L_20_5,
    output F2Adef_L_20_6,
    output F2Adef_L_21_0,
    output F2Adef_L_21_1,
    output F2Adef_L_21_2,
    output F2Adef_L_21_3,
    output F2Adef_L_22_0,
    output F2Adef_L_22_1,
    output F2Adef_L_22_2,
    output F2Adef_L_22_3,
    output F2Adef_L_22_4,
    output F2Adef_L_22_5,
    output F2Adef_L_22_6,
    output F2Adef_L_23_0,
    output F2Adef_L_23_1,
    output F2Adef_L_23_2,
    output F2Adef_L_23_3,
    output F2Adef_L_24_0,
    output F2Adef_L_24_1,
    output F2Adef_L_24_2,
    output F2Adef_L_24_3,
    output F2Adef_L_24_4,
    output F2Adef_L_24_5,
    output F2Adef_L_24_6,
    output F2Adef_L_25_0,
    output F2Adef_L_25_1,
    output F2Adef_L_25_2,
    output F2Adef_L_25_3,
    output F2Adef_L_26_0,
    output F2Adef_L_26_1,
    output F2Adef_L_26_2,
    output F2Adef_L_26_3,
    output F2Adef_L_26_4,
    output F2Adef_L_26_5,
    output F2Adef_L_26_6,
    output F2Adef_L_27_0,
    output F2Adef_L_27_1,
    output F2Adef_L_27_2,
    output F2Adef_L_27_3,
    output F2Adef_L_28_0,
    output F2Adef_L_28_1,
    output F2Adef_L_28_2,
    output F2Adef_L_28_3,
    output F2Adef_L_28_4,
    output F2Adef_L_28_5,
    output F2Adef_L_28_6,
    output F2Adef_L_29_0,
    output F2Adef_L_29_1,
    output F2Adef_L_29_2,
    output F2Adef_L_29_3,
    output F2Adef_L_2_0,
    output F2Adef_L_2_1,
    output F2Adef_L_2_2,
    output F2Adef_L_2_3,
    output F2Adef_L_2_4,
    output F2Adef_L_2_5,
    output F2Adef_L_2_6,
    output F2Adef_L_30_0,
    output F2Adef_L_30_1,
    output F2Adef_L_30_2,
    output F2Adef_L_30_3,
    output F2Adef_L_30_4,
    output F2Adef_L_30_5,
    output F2Adef_L_30_6,
    output F2Adef_L_31_0,
    output F2Adef_L_31_1,
    output F2Adef_L_31_2,
    output F2Adef_L_31_3,
    output F2Adef_L_32_0,
    output F2Adef_L_32_1,
    output F2Adef_L_32_2,
    output F2Adef_L_32_3,
    output F2Adef_L_32_4,
    output F2Adef_L_32_5,
    output F2Adef_L_32_6,
    output F2Adef_L_3_0,
    output F2Adef_L_3_1,
    output F2Adef_L_3_2,
    output F2Adef_L_3_3,
    output F2Adef_L_4_0,
    output F2Adef_L_4_1,
    output F2Adef_L_4_2,
    output F2Adef_L_4_3,
    output F2Adef_L_4_4,
    output F2Adef_L_4_5,
    output F2Adef_L_4_6,
    output F2Adef_L_5_0,
    output F2Adef_L_5_1,
    output F2Adef_L_5_2,
    output F2Adef_L_5_3,
    output F2Adef_L_6_0,
    output F2Adef_L_6_1,
    output F2Adef_L_6_2,
    output F2Adef_L_6_3,
    output F2Adef_L_6_4,
    output F2Adef_L_6_5,
    output F2Adef_L_6_6,
    output F2Adef_L_7_0,
    output F2Adef_L_7_1,
    output F2Adef_L_7_2,
    output F2Adef_L_7_3,
    output F2Adef_L_8_0,
    output F2Adef_L_8_1,
    output F2Adef_L_8_2,
    output F2Adef_L_8_3,
    output F2Adef_L_8_4,
    output F2Adef_L_8_5,
    output F2Adef_L_8_6,
    output F2Adef_L_9_0,
    output F2Adef_L_9_1,
    output F2Adef_L_9_2,
    output F2Adef_L_9_3,
    output F2Adef_R_10_0,
    output F2Adef_R_10_1,
    output F2Adef_R_10_2,
    output F2Adef_R_10_3,
    output F2Adef_R_10_4,
    output F2Adef_R_10_5,
    output F2Adef_R_10_6,
    output F2Adef_R_11_0,
    output F2Adef_R_11_1,
    output F2Adef_R_11_2,
    output F2Adef_R_11_3,
    output F2Adef_R_12_0,
    output F2Adef_R_12_1,
    output F2Adef_R_12_2,
    output F2Adef_R_12_3,
    output F2Adef_R_12_4,
    output F2Adef_R_12_5,
    output F2Adef_R_12_6,
    output F2Adef_R_13_0,
    output F2Adef_R_13_1,
    output F2Adef_R_13_2,
    output F2Adef_R_13_3,
    output F2Adef_R_14_0,
    output F2Adef_R_14_1,
    output F2Adef_R_14_2,
    output F2Adef_R_14_3,
    output F2Adef_R_14_4,
    output F2Adef_R_14_5,
    output F2Adef_R_14_6,
    output F2Adef_R_15_0,
    output F2Adef_R_15_1,
    output F2Adef_R_15_2,
    output F2Adef_R_15_3,
    output F2Adef_R_16_0,
    output F2Adef_R_16_1,
    output F2Adef_R_16_2,
    output F2Adef_R_16_3,
    output F2Adef_R_16_4,
    output F2Adef_R_16_5,
    output F2Adef_R_16_6,
    output F2Adef_R_17_0,
    output F2Adef_R_17_1,
    output F2Adef_R_17_2,
    output F2Adef_R_17_3,
    output F2Adef_R_18_0,
    output F2Adef_R_18_1,
    output F2Adef_R_18_2,
    output F2Adef_R_18_3,
    output F2Adef_R_18_4,
    output F2Adef_R_18_5,
    output F2Adef_R_18_6,
    output F2Adef_R_19_0,
    output F2Adef_R_19_1,
    output F2Adef_R_19_2,
    output F2Adef_R_19_3,
    output F2Adef_R_1_0,
    output F2Adef_R_1_1,
    output F2Adef_R_1_2,
    output F2Adef_R_1_3,
    output F2Adef_R_20_0,
    output F2Adef_R_20_1,
    output F2Adef_R_20_2,
    output F2Adef_R_20_3,
    output F2Adef_R_20_4,
    output F2Adef_R_20_5,
    output F2Adef_R_20_6,
    output F2Adef_R_21_0,
    output F2Adef_R_21_1,
    output F2Adef_R_21_2,
    output F2Adef_R_21_3,
    output F2Adef_R_22_0,
    output F2Adef_R_22_1,
    output F2Adef_R_22_2,
    output F2Adef_R_22_3,
    output F2Adef_R_22_4,
    output F2Adef_R_22_5,
    output F2Adef_R_22_6,
    output F2Adef_R_23_0,
    output F2Adef_R_23_1,
    output F2Adef_R_23_2,
    output F2Adef_R_23_3,
    output F2Adef_R_24_0,
    output F2Adef_R_24_1,
    output F2Adef_R_24_2,
    output F2Adef_R_24_3,
    output F2Adef_R_24_4,
    output F2Adef_R_24_5,
    output F2Adef_R_24_6,
    output F2Adef_R_25_0,
    output F2Adef_R_25_1,
    output F2Adef_R_25_2,
    output F2Adef_R_25_3,
    output F2Adef_R_26_0,
    output F2Adef_R_26_1,
    output F2Adef_R_26_2,
    output F2Adef_R_26_3,
    output F2Adef_R_26_4,
    output F2Adef_R_26_5,
    output F2Adef_R_26_6,
    output F2Adef_R_27_0,
    output F2Adef_R_27_1,
    output F2Adef_R_27_2,
    output F2Adef_R_27_3,
    output F2Adef_R_28_0,
    output F2Adef_R_28_1,
    output F2Adef_R_28_2,
    output F2Adef_R_28_3,
    output F2Adef_R_28_4,
    output F2Adef_R_28_5,
    output F2Adef_R_28_6,
    output F2Adef_R_29_0,
    output F2Adef_R_29_1,
    output F2Adef_R_29_2,
    output F2Adef_R_29_3,
    output F2Adef_R_2_0,
    output F2Adef_R_2_1,
    output F2Adef_R_2_2,
    output F2Adef_R_2_3,
    output F2Adef_R_2_4,
    output F2Adef_R_2_5,
    output F2Adef_R_2_6,
    output F2Adef_R_30_0,
    output F2Adef_R_30_1,
    output F2Adef_R_30_2,
    output F2Adef_R_30_3,
    output F2Adef_R_30_4,
    output F2Adef_R_30_5,
    output F2Adef_R_30_6,
    output F2Adef_R_31_0,
    output F2Adef_R_31_1,
    output F2Adef_R_31_2,
    output F2Adef_R_31_3,
    output F2Adef_R_32_0,
    output F2Adef_R_32_1,
    output F2Adef_R_32_2,
    output F2Adef_R_32_3,
    output F2Adef_R_32_4,
    output F2Adef_R_32_5,
    output F2Adef_R_32_6,
    output F2Adef_R_3_0,
    output F2Adef_R_3_1,
    output F2Adef_R_3_2,
    output F2Adef_R_3_3,
    output F2Adef_R_4_0,
    output F2Adef_R_4_1,
    output F2Adef_R_4_2,
    output F2Adef_R_4_3,
    output F2Adef_R_4_4,
    output F2Adef_R_4_5,
    output F2Adef_R_4_6,
    output F2Adef_R_5_0,
    output F2Adef_R_5_1,
    output F2Adef_R_5_2,
    output F2Adef_R_5_3,
    output F2Adef_R_6_0,
    output F2Adef_R_6_1,
    output F2Adef_R_6_2,
    output F2Adef_R_6_3,
    output F2Adef_R_6_4,
    output F2Adef_R_6_5,
    output F2Adef_R_6_6,
    output F2Adef_R_7_0,
    output F2Adef_R_7_1,
    output F2Adef_R_7_2,
    output F2Adef_R_7_3,
    output F2Adef_R_8_0,
    output F2Adef_R_8_1,
    output F2Adef_R_8_2,
    output F2Adef_R_8_3,
    output F2Adef_R_8_4,
    output F2Adef_R_8_5,
    output F2Adef_R_8_6,
    output F2Adef_R_9_0,
    output F2Adef_R_9_1,
    output F2Adef_R_9_2,
    output F2Adef_R_9_3,
    output F2Adef_T_10_0,
    output F2Adef_T_10_1,
    output F2Adef_T_10_2,
    output F2Adef_T_10_3,
    output F2Adef_T_10_4,
    output F2Adef_T_10_5,
    output F2Adef_T_10_6,
    output F2Adef_T_11_0,
    output F2Adef_T_11_1,
    output F2Adef_T_11_2,
    output F2Adef_T_11_3,
    output F2Adef_T_12_0,
    output F2Adef_T_12_1,
    output F2Adef_T_12_2,
    output F2Adef_T_12_3,
    output F2Adef_T_12_4,
    output F2Adef_T_12_5,
    output F2Adef_T_12_6,
    output F2Adef_T_13_0,
    output F2Adef_T_13_1,
    output F2Adef_T_13_2,
    output F2Adef_T_13_3,
    output F2Adef_T_14_0,
    output F2Adef_T_14_1,
    output F2Adef_T_14_2,
    output F2Adef_T_14_3,
    output F2Adef_T_14_4,
    output F2Adef_T_14_5,
    output F2Adef_T_14_6,
    output F2Adef_T_15_0,
    output F2Adef_T_15_1,
    output F2Adef_T_15_2,
    output F2Adef_T_15_3,
    output F2Adef_T_16_0,
    output F2Adef_T_16_1,
    output F2Adef_T_16_2,
    output F2Adef_T_16_3,
    output F2Adef_T_16_4,
    output F2Adef_T_16_5,
    output F2Adef_T_16_6,
    output F2Adef_T_17_0,
    output F2Adef_T_17_1,
    output F2Adef_T_17_2,
    output F2Adef_T_17_3,
    output F2Adef_T_18_0,
    output F2Adef_T_18_1,
    output F2Adef_T_18_2,
    output F2Adef_T_18_3,
    output F2Adef_T_18_4,
    output F2Adef_T_18_5,
    output F2Adef_T_18_6,
    output F2Adef_T_19_0,
    output F2Adef_T_19_1,
    output F2Adef_T_19_2,
    output F2Adef_T_19_3,
    output F2Adef_T_1_0,
    output F2Adef_T_1_1,
    output F2Adef_T_1_2,
    output F2Adef_T_1_3,
    output F2Adef_T_20_0,
    output F2Adef_T_20_1,
    output F2Adef_T_20_2,
    output F2Adef_T_20_3,
    output F2Adef_T_20_4,
    output F2Adef_T_20_5,
    output F2Adef_T_20_6,
    output F2Adef_T_21_0,
    output F2Adef_T_21_1,
    output F2Adef_T_21_2,
    output F2Adef_T_21_3,
    output F2Adef_T_22_0,
    output F2Adef_T_22_1,
    output F2Adef_T_22_2,
    output F2Adef_T_22_3,
    output F2Adef_T_22_4,
    output F2Adef_T_22_5,
    output F2Adef_T_22_6,
    output F2Adef_T_23_0,
    output F2Adef_T_23_1,
    output F2Adef_T_23_2,
    output F2Adef_T_23_3,
    output F2Adef_T_24_0,
    output F2Adef_T_24_1,
    output F2Adef_T_24_2,
    output F2Adef_T_24_3,
    output F2Adef_T_24_4,
    output F2Adef_T_24_5,
    output F2Adef_T_24_6,
    output F2Adef_T_25_0,
    output F2Adef_T_25_1,
    output F2Adef_T_25_2,
    output F2Adef_T_25_3,
    output F2Adef_T_26_0,
    output F2Adef_T_26_1,
    output F2Adef_T_26_2,
    output F2Adef_T_26_3,
    output F2Adef_T_26_4,
    output F2Adef_T_26_5,
    output F2Adef_T_26_6,
    output F2Adef_T_27_0,
    output F2Adef_T_27_1,
    output F2Adef_T_27_2,
    output F2Adef_T_27_3,
    output F2Adef_T_28_0,
    output F2Adef_T_28_1,
    output F2Adef_T_28_2,
    output F2Adef_T_28_3,
    output F2Adef_T_28_4,
    output F2Adef_T_28_5,
    output F2Adef_T_28_6,
    output F2Adef_T_29_0,
    output F2Adef_T_29_1,
    output F2Adef_T_29_2,
    output F2Adef_T_29_3,
    output F2Adef_T_2_0,
    output F2Adef_T_2_1,
    output F2Adef_T_2_2,
    output F2Adef_T_2_3,
    output F2Adef_T_2_4,
    output F2Adef_T_2_5,
    output F2Adef_T_2_6,
    output F2Adef_T_30_0,
    output F2Adef_T_30_1,
    output F2Adef_T_30_2,
    output F2Adef_T_30_3,
    output F2Adef_T_30_4,
    output F2Adef_T_30_5,
    output F2Adef_T_30_6,
    output F2Adef_T_31_0,
    output F2Adef_T_31_1,
    output F2Adef_T_31_2,
    output F2Adef_T_31_3,
    output F2Adef_T_32_0,
    output F2Adef_T_32_1,
    output F2Adef_T_32_2,
    output F2Adef_T_32_3,
    output F2Adef_T_32_4,
    output F2Adef_T_32_5,
    output F2Adef_T_32_6,
    output F2Adef_T_3_0,
    output F2Adef_T_3_1,
    output F2Adef_T_3_2,
    output F2Adef_T_3_3,
    output F2Adef_T_4_0,
    output F2Adef_T_4_1,
    output F2Adef_T_4_2,
    output F2Adef_T_4_3,
    output F2Adef_T_4_4,
    output F2Adef_T_4_5,
    output F2Adef_T_4_6,
    output F2Adef_T_5_0,
    output F2Adef_T_5_1,
    output F2Adef_T_5_2,
    output F2Adef_T_5_3,
    output F2Adef_T_6_0,
    output F2Adef_T_6_1,
    output F2Adef_T_6_2,
    output F2Adef_T_6_3,
    output F2Adef_T_6_4,
    output F2Adef_T_6_5,
    output F2Adef_T_6_6,
    output F2Adef_T_7_0,
    output F2Adef_T_7_1,
    output F2Adef_T_7_2,
    output F2Adef_T_7_3,
    output F2Adef_T_8_0,
    output F2Adef_T_8_1,
    output F2Adef_T_8_2,
    output F2Adef_T_8_3,
    output F2Adef_T_8_4,
    output F2Adef_T_8_5,
    output F2Adef_T_8_6,
    output F2Adef_T_9_0,
    output F2Adef_T_9_1,
    output F2Adef_T_9_2,
    output F2Adef_T_9_3,
    output F2Areg_B_11_0,
    output F2Areg_B_11_1,
    output F2Areg_B_13_0,
    output F2Areg_B_13_1,
    output F2Areg_B_15_0,
    output F2Areg_B_15_1,
    output F2Areg_B_17_0,
    output F2Areg_B_17_1,
    output F2Areg_B_19_0,
    output F2Areg_B_19_1,
    output F2Areg_B_1_0,
    output F2Areg_B_1_1,
    output F2Areg_B_21_0,
    output F2Areg_B_21_1,
    output F2Areg_B_23_0,
    output F2Areg_B_23_1,
    output F2Areg_B_25_0,
    output F2Areg_B_25_1,
    output F2Areg_B_27_0,
    output F2Areg_B_27_1,
    output F2Areg_B_29_0,
    output F2Areg_B_29_1,
    output F2Areg_B_31_0,
    output F2Areg_B_31_1,
    output F2Areg_B_3_0,
    output F2Areg_B_3_1,
    output F2Areg_B_5_0,
    output F2Areg_B_5_1,
    output F2Areg_B_7_0,
    output F2Areg_B_7_1,
    output F2Areg_B_9_0,
    output F2Areg_B_9_1,
    output F2Areg_L_11_0,
    output F2Areg_L_11_1,
    output F2Areg_L_13_0,
    output F2Areg_L_13_1,
    output F2Areg_L_15_0,
    output F2Areg_L_15_1,
    output F2Areg_L_17_0,
    output F2Areg_L_17_1,
    output F2Areg_L_19_0,
    output F2Areg_L_19_1,
    output F2Areg_L_1_0,
    output F2Areg_L_1_1,
    output F2Areg_L_21_0,
    output F2Areg_L_21_1,
    output F2Areg_L_23_0,
    output F2Areg_L_23_1,
    output F2Areg_L_25_0,
    output F2Areg_L_25_1,
    output F2Areg_L_27_0,
    output F2Areg_L_27_1,
    output F2Areg_L_29_0,
    output F2Areg_L_29_1,
    output F2Areg_L_31_0,
    output F2Areg_L_31_1,
    output F2Areg_L_3_0,
    output F2Areg_L_3_1,
    output F2Areg_L_5_0,
    output F2Areg_L_5_1,
    output F2Areg_L_7_0,
    output F2Areg_L_7_1,
    output F2Areg_L_9_0,
    output F2Areg_L_9_1,
    output F2Areg_R_11_0,
    output F2Areg_R_11_1,
    output F2Areg_R_13_0,
    output F2Areg_R_13_1,
    output F2Areg_R_15_0,
    output F2Areg_R_15_1,
    output F2Areg_R_17_0,
    output F2Areg_R_17_1,
    output F2Areg_R_19_0,
    output F2Areg_R_19_1,
    output F2Areg_R_1_0,
    output F2Areg_R_1_1,
    output F2Areg_R_21_0,
    output F2Areg_R_21_1,
    output F2Areg_R_23_0,
    output F2Areg_R_23_1,
    output F2Areg_R_25_0,
    output F2Areg_R_25_1,
    output F2Areg_R_27_0,
    output F2Areg_R_27_1,
    output F2Areg_R_29_0,
    output F2Areg_R_29_1,
    output F2Areg_R_31_0,
    output F2Areg_R_31_1,
    output F2Areg_R_3_0,
    output F2Areg_R_3_1,
    output F2Areg_R_5_0,
    output F2Areg_R_5_1,
    output F2Areg_R_7_0,
    output F2Areg_R_7_1,
    output F2Areg_R_9_0,
    output F2Areg_R_9_1,
    output F2Areg_T_11_0,
    output F2Areg_T_11_1,
    output F2Areg_T_13_0,
    output F2Areg_T_13_1,
    output F2Areg_T_15_0,
    output F2Areg_T_15_1,
    output F2Areg_T_17_0,
    output F2Areg_T_17_1,
    output F2Areg_T_19_0,
    output F2Areg_T_19_1,
    output F2Areg_T_1_0,
    output F2Areg_T_1_1,
    output F2Areg_T_21_0,
    output F2Areg_T_21_1,
    output F2Areg_T_23_0,
    output F2Areg_T_23_1,
    output F2Areg_T_25_0,
    output F2Areg_T_25_1,
    output F2Areg_T_27_0,
    output F2Areg_T_27_1,
    output F2Areg_T_29_0,
    output F2Areg_T_29_1,
    output F2Areg_T_31_0,
    output F2Areg_T_31_1,
    output F2Areg_T_3_0,
    output F2Areg_T_3_1,
    output F2Areg_T_5_0,
    output F2Areg_T_5_1,
    output F2Areg_T_7_0,
    output F2Areg_T_7_1,
    output F2Areg_T_9_0,
    output F2Areg_T_9_1,
    output BL_DOUT_0_,
    output BL_DOUT_1_,
    output BL_DOUT_2_,
    output BL_DOUT_3_,
    output BL_DOUT_4_,
    output BL_DOUT_5_,
    output BL_DOUT_6_,
    output BL_DOUT_7_,
    output BL_DOUT_8_,
    output BL_DOUT_9_,
    output BL_DOUT_10_,
    output BL_DOUT_11_,
    output BL_DOUT_12_,
    output BL_DOUT_13_,
    output BL_DOUT_14_,
    output BL_DOUT_15_,
    output BL_DOUT_16_,
    output BL_DOUT_17_,
    output BL_DOUT_18_,
    output BL_DOUT_19_,
    output BL_DOUT_20_,
    output BL_DOUT_21_,
    output BL_DOUT_22_,
    output BL_DOUT_23_,
    output BL_DOUT_24_,
    output BL_DOUT_25_,
    output BL_DOUT_26_,
    output BL_DOUT_27_,
    output BL_DOUT_28_,
    output BL_DOUT_29_,
    output BL_DOUT_30_,
    output BL_DOUT_31_,
    output FB_SPE_OUT_0_,
    output FB_SPE_OUT_1_,
    output FB_SPE_OUT_2_,
    output FB_SPE_OUT_3_,
    output PARALLEL_CFG,
    input  BL_CLK,
    input  BL_DIN_0_,
    input  BL_DIN_1_,
    input  BL_DIN_2_,
    input  BL_DIN_3_,
    input  BL_DIN_4_,
    input  BL_DIN_5_,
    input  BL_DIN_6_,
    input  BL_DIN_7_,
    input  BL_DIN_8_,
    input  BL_DIN_9_,
    input  BL_DIN_10_,
    input  BL_DIN_11_,
    input  BL_DIN_12_,
    input  BL_DIN_13_,
    input  BL_DIN_14_,
    input  BL_DIN_15_,
    input  BL_DIN_16_,
    input  BL_DIN_17_,
    input  BL_DIN_18_,
    input  BL_DIN_19_,
    input  BL_DIN_20_,
    input  BL_DIN_21_,
    input  BL_DIN_22_,
    input  BL_DIN_23_,
    input  BL_DIN_24_,
    input  BL_DIN_25_,
    input  BL_DIN_26_,
    input  BL_DIN_27_,
    input  BL_DIN_28_,
    input  BL_DIN_29_,
    input  BL_DIN_30_,
    input  BL_DIN_31_,
    input  BL_PWRGATE_0_,
    input  BL_PWRGATE_1_,
    input  BL_PWRGATE_2_,
    input  BL_PWRGATE_3_,
    input  CLOAD_DIN_SEL,
    input  DIN_INT_L_ONLY,
    input  DIN_INT_R_ONLY,
    input  DIN_SLC_TB_INT,
    input  FB_CFG_DONE,
    input  FB_ISO_ENB,
    input  FB_SPE_IN_0_,
    input  FB_SPE_IN_1_,
    input  FB_SPE_IN_2_,
    input  FB_SPE_IN_3_,
    input  ISO_EN_0_,
    input  ISO_EN_1_,
    input  ISO_EN_2_,
    input  ISO_EN_3_,
    input  M_0_,
    input  M_1_,
    input  M_2_,
    input  M_3_,
    input  M_4_,
    input  M_5_,
    input  MLATCH,
    input  PB,
    input  NB,
    input  PCHG_B,
    input  PI_PWR_0_,
    input  PI_PWR_1_,
    input  PI_PWR_2_,
    input  PI_PWR_3_,
    input  POR,
    input  PROG_0_,
    input  PROG_1_,
    input  PROG_2_,
    input  PROG_3_,
    input  PROG_IFX,
    input  PWR_GATE,
    input  RE,
    input  STM,
    input  VLP_CLKDIS_0_,
    input  VLP_CLKDIS_1_,
    input  VLP_CLKDIS_2_,
    input  VLP_CLKDIS_3_,
    input  VLP_CLKDIS_IFX,
    input  VLP_PWRDIS_0_,
    input  VLP_PWRDIS_1_,
    input  VLP_PWRDIS_2_,
    input  VLP_PWRDIS_3_,
    input  VLP_PWRDIS_IFX,
    input  VLP_SRDIS_0_,
    input  VLP_SRDIS_1_,
    input  VLP_SRDIS_2_,
    input  VLP_SRDIS_3_,
    input  VLP_SRDIS_IFX,
    input  WE,
    input  WE_INT,
    input  WL_CLK,
    input  WL_CLOAD_SEL_0_,
    input  WL_CLOAD_SEL_1_,
    input  WL_CLOAD_SEL_2_,
    input  WL_DIN_0_,
    input  WL_DIN_1_,
    input  WL_DIN_2_,
    input  WL_DIN_3_,
    input  WL_DIN_4_,
    input  WL_DIN_5_,
    input  WL_EN,
    input  WL_INT_DIN_SEL,
    input  WL_PWRGATE_0_,
    input  WL_PWRGATE_1_,
    input  WL_RESETB,
    input  WL_SEL_0_,
    input  WL_SEL_1_,
    input  WL_SEL_2_,
    input  WL_SEL_3_,
    input  WL_SEL_TB_INT
);


  top top1_rtl (
      //	top1 top1_vq (
      .RESET({A2F_L_2_4, A2F_L_25_2, A2F_R_29_2, A2F_R_6_0}),
      .lint_GNT(F2A_L_15_8),
      .lint_REQ(A2F_L_12_2),
      .lint_VALID(F2A_L_14_9),
      .lint_WEN(A2F_L_12_3),
      .lint_clk(F2A_L_14_0),
      .m0_coef_powerdn(F2Adef_T_13_0),
      .m0_coef_rclk(F2A_T_15_0),
      .m0_coef_wclk(F2A_T_13_0),
      .m0_coef_wdsel(F2A_T_14_11),
      .m0_coef_we(F2A_T_14_10),
      .m0_m0_clk(F2A_T_7_0),
      .m0_m0_clken(F2A_T_6_5),
      .m0_m0_clr(F2A_T_6_14),
      .m0_m0_csel(F2A_T_9_0),
      .m0_m0_osel(F2A_T_6_4),
      .m0_m0_reset(F2A_T_11_6),
      .m0_m0_rnd(F2A_T_6_13),
      .m0_m0_sat(F2A_T_6_12),
      .m0_m0_tc(F2A_T_11_5),
      .m0_m1_clk(F2A_T_19_0),
      .m0_m1_clken(F2A_T_18_17),
      .m0_m1_clr(F2A_T_18_16),
      .m0_m1_csel(F2A_T_21_7),
      .m0_m1_osel(F2A_T_19_1),
      .m0_m1_reset(F2A_T_19_3),
      .m0_m1_rnd(F2A_T_18_15),
      .m0_m1_sat(F2A_T_18_14),
      .m0_m1_tc(F2A_T_19_2),
      .m0_oper0_powerdn(F2Adef_T_6_1),
      .m0_oper0_rclk(F2A_T_6_0),
      .m0_oper0_wclk(F2A_T_2_0),
      .m0_oper0_wdsel(F2A_T_2_3),
      .m0_oper0_we(F2A_T_5_2),
      .m0_oper1_powerdn(F2Adef_T_24_0),
      .m0_oper1_rclk(F2A_T_29_0),
      .m0_oper1_wclk(F2A_T_28_0),
      .m0_oper1_wdsel(F2A_T_28_3),
      .m0_oper1_we(F2A_T_28_4),
      .m1_coef_powerdn(F2Adef_B_13_0),
      .m1_coef_rclk(F2A_B_15_0),
      .m1_coef_wclk(F2A_B_13_0),
      .m1_coef_wdsel(F2A_B_14_11),
      .m1_coef_we(F2A_B_14_10),
      .m1_m0_clk(F2A_B_7_0),
      .m1_m0_clken(F2A_B_6_5),
      .m1_m0_clr(F2A_B_6_14),
      .m1_m0_csel(F2A_B_9_0),
      .m1_m0_osel(F2A_B_6_4),
      .m1_m0_reset(F2A_B_11_6),
      .m1_m0_rnd(F2A_B_6_13),
      .m1_m0_sat(F2A_B_6_12),
      .m1_m0_tc(F2A_B_11_5),
      .m1_m1_clk(F2A_B_19_0),
      .m1_m1_clken(F2A_B_18_16),
      .m1_m1_clr(F2A_B_18_15),
      .m1_m1_csel(F2A_B_21_7),
      .m1_m1_osel(F2A_B_19_1),
      .m1_m1_reset(F2A_B_19_3),
      .m1_m1_rnd(F2A_B_18_14),
      .m1_m1_sat(F2A_B_18_13),
      .m1_m1_tc(F2A_B_19_2),
      .m1_oper0_powerdn(F2Adef_B_6_1),
      .m1_oper0_rclk(F2A_B_6_0),
      .m1_oper0_wclk(F2A_B_2_0),
      .m1_oper0_wdsel(F2A_B_2_3),
      .m1_oper0_we(F2A_B_5_2),
      .m1_oper1_powerdn(F2Adef_B_24_1),
      .m1_oper1_rclk(F2A_B_29_0),
      .m1_oper1_wclk(F2A_B_28_0),
      .m1_oper1_wdsel(F2A_B_28_3),
      .m1_oper1_we(F2A_B_28_4),
      .tcdm_clk_p0(F2A_R_3_0),
      .tcdm_clk_p1(F2A_R_9_0),
      .tcdm_clk_p2(F2A_R_17_0),
      .tcdm_clk_p3(F2A_R_23_0),
      .tcdm_gnt_p0(A2F_R_3_5),
      .tcdm_gnt_p1(A2F_R_9_5),
      .tcdm_gnt_p2(A2F_R_17_5),
      .tcdm_gnt_p3(A2F_R_23_5),
      .tcdm_req_p0(F2A_R_3_1),
      .tcdm_req_p1(F2A_R_9_1),
      .tcdm_req_p2(F2A_R_17_1),
      .tcdm_req_p3(F2A_R_23_1),
      .tcdm_valid_p0(A2F_R_3_4),
      .tcdm_valid_p1(A2F_R_9_4),
      .tcdm_valid_p2(A2F_R_17_4),
      .tcdm_valid_p3(A2F_R_23_4),
      .tcdm_wen_p0(F2A_R_3_2),
      .tcdm_wen_p1(F2A_R_9_2),
      .tcdm_wen_p2(F2A_R_17_2),
      .tcdm_wen_p3(F2A_R_23_2),
      .tcdm_fmo_p0(A2F_R_5_4),
      .tcdm_fmo_p1(A2F_R_11_4),
      .tcdm_fmo_p2(A2F_R_19_4),
      .tcdm_fmo_p3(A2F_R_25_4),
      .CLK({A2F_CLK5, A2F_CLK4, A2F_CLK3, A2F_CLK2, A2F_CLK1, A2F_CLK0}),
      .control_in({
        A2F_L_23_4,
        A2F_L_23_3,
        A2F_L_23_2,
        A2F_L_23_1,
        A2F_L_23_0,
        A2F_L_22_6,
        A2F_L_22_5,
        A2F_L_22_4,
        A2F_L_22_3,
        A2F_L_22_2,
        A2F_L_22_1,
        A2F_L_22_0,
        A2F_L_21_5,
        A2F_L_21_4,
        A2F_L_21_3,
        A2F_L_21_2,
        A2F_L_21_1,
        A2F_L_21_0,
        A2F_L_20_7,
        A2F_L_20_6,
        A2F_L_20_5,
        A2F_L_20_4,
        A2F_L_20_3,
        A2F_L_20_2,
        A2F_L_20_1,
        A2F_L_20_0,
        A2F_L_19_5,
        A2F_L_19_4,
        A2F_L_19_3,
        A2F_L_19_2,
        A2F_L_19_1,
        A2F_L_19_0
      }),
      .events_o({
        F2A_L_32_8,
        F2A_L_31_8,
        F2A_L_30_8,
        F2A_L_29_8,
        F2A_L_28_8,
        F2A_L_27_8,
        F2A_L_26_8,
        F2A_L_25_8,
        F2A_L_8_8,
        F2A_L_6_17,
        F2A_L_6_8,
        F2A_L_5_11,
        F2A_L_5_2,
        F2A_L_4_8,
        F2A_L_3_8,
        F2A_L_2_8
      }),
      .fpgaio_in({
        A2F_L_18_1,
        A2F_L_18_0,
        A2F_L_17_5,
        A2F_L_17_4,
        A2F_L_17_3,
        A2F_L_17_2,
        A2F_L_17_1,
        A2F_L_17_0,
        A2F_L_16_7,
        A2F_L_16_6,
        A2F_L_16_5,
        A2F_L_16_4,
        A2F_L_16_3,
        A2F_L_16_2,
        A2F_L_16_1,
        A2F_L_16_0,
        A2F_L_32_3,
        A2F_L_32_2,
        A2F_L_32_1,
        A2F_L_32_0,
        A2F_L_31_3,
        A2F_L_31_2,
        A2F_L_31_1,
        A2F_L_31_0,
        A2F_L_30_3,
        A2F_L_30_2,
        A2F_L_30_1,
        A2F_L_30_0,
        A2F_L_29_3,
        A2F_L_29_2,
        A2F_L_29_1,
        A2F_L_29_0,
        A2F_L_28_3,
        A2F_L_28_2,
        A2F_L_28_1,
        A2F_L_28_0,
        A2F_L_27_3,
        A2F_L_27_2,
        A2F_L_27_1,
        A2F_L_27_0,
        A2F_L_26_3,
        A2F_L_26_2,
        A2F_L_26_1,
        A2F_L_26_0,
        A2F_L_25_4,
        A2F_L_25_3,
        A2F_L_25_1,
        A2F_L_25_0,
        A2F_L_7_3,
        A2F_L_7_2,
        A2F_L_7_1,
        A2F_L_7_0,
        A2F_L_6_5,
        A2F_L_6_4,
        A2F_L_6_3,
        A2F_L_6_2,
        A2F_L_6_1,
        A2F_L_6_0,
        A2F_L_5_5,
        A2F_L_5_4,
        A2F_L_5_3,
        A2F_L_5_2,
        A2F_L_5_1,
        A2F_L_5_0,
        A2F_L_4_7,
        A2F_L_4_6,
        A2F_L_4_5,
        A2F_L_4_4,
        A2F_L_4_3,
        A2F_L_4_2,
        A2F_L_3_5,
        A2F_L_3_4,
        A2F_L_3_3,
        A2F_L_3_2,
        A2F_L_3_1,
        A2F_L_3_0,
        A2F_L_2_3,
        A2F_L_2_2,
        A2F_L_2_1,
        A2F_L_2_0
      }),
      .fpgaio_oe({
        F2A_L_19_7,
        F2A_L_19_5,
        F2A_L_19_3,
        F2A_L_19_1,
        F2A_L_18_15,
        F2A_L_18_13,
        F2A_L_18_11,
        F2A_L_18_9,
        F2A_L_18_7,
        F2A_L_18_5,
        F2A_L_18_3,
        F2A_L_18_1,
        F2A_L_17_7,
        F2A_L_17_5,
        F2A_L_17_3,
        F2A_L_17_1,
        F2A_L_32_7,
        F2A_L_32_5,
        F2A_L_32_3,
        F2A_L_32_1,
        F2A_L_31_7,
        F2A_L_31_5,
        F2A_L_31_3,
        F2A_L_31_1,
        F2A_L_30_7,
        F2A_L_30_5,
        F2A_L_30_3,
        F2A_L_30_1,
        F2A_L_29_7,
        F2A_L_29_5,
        F2A_L_29_3,
        F2A_L_29_1,
        F2A_L_28_7,
        F2A_L_28_5,
        F2A_L_28_3,
        F2A_L_28_1,
        F2A_L_27_7,
        F2A_L_27_5,
        F2A_L_27_3,
        F2A_L_27_1,
        F2A_L_26_7,
        F2A_L_26_5,
        F2A_L_26_3,
        F2A_L_26_1,
        F2A_L_25_7,
        F2A_L_25_5,
        F2A_L_25_3,
        F2A_L_25_1,
        F2A_L_8_7,
        F2A_L_8_5,
        F2A_L_8_3,
        F2A_L_8_1,
        F2A_L_6_16,
        F2A_L_6_14,
        F2A_L_6_12,
        F2A_L_6_10,
        F2A_L_6_7,
        F2A_L_6_5,
        F2A_L_6_3,
        F2A_L_6_1,
        F2A_L_5_10,
        F2A_L_5_8,
        F2A_L_5_6,
        F2A_L_5_4,
        F2A_L_5_1,
        F2A_L_4_14,
        F2A_L_4_12,
        F2A_L_4_10,
        F2A_L_4_7,
        F2A_L_4_5,
        F2A_L_4_3,
        F2A_L_4_1,
        F2A_L_3_7,
        F2A_L_3_5,
        F2A_L_3_3,
        F2A_L_3_1,
        F2A_L_2_7,
        F2A_L_2_5,
        F2A_L_2_3,
        F2A_L_2_1
      }),
      .fpgaio_out({
        F2A_L_19_6,
        F2A_L_19_4,
        F2A_L_19_2,
        F2A_L_19_0,
        F2A_L_18_14,
        F2A_L_18_12,
        F2A_L_18_10,
        F2A_L_18_8,
        F2A_L_18_6,
        F2A_L_18_4,
        F2A_L_18_2,
        F2A_L_18_0,
        F2A_L_17_6,
        F2A_L_17_4,
        F2A_L_17_2,
        F2A_L_17_0,
        F2A_L_32_6,
        F2A_L_32_4,
        F2A_L_32_2,
        F2A_L_32_0,
        F2A_L_31_6,
        F2A_L_31_4,
        F2A_L_31_2,
        F2A_L_31_0,
        F2A_L_30_6,
        F2A_L_30_4,
        F2A_L_30_2,
        F2A_L_30_0,
        F2A_L_29_6,
        F2A_L_29_4,
        F2A_L_29_2,
        F2A_L_29_0,
        F2A_L_28_6,
        F2A_L_28_4,
        F2A_L_28_2,
        F2A_L_28_0,
        F2A_L_27_6,
        F2A_L_27_4,
        F2A_L_27_2,
        F2A_L_27_0,
        F2A_L_26_6,
        F2A_L_26_4,
        F2A_L_26_2,
        F2A_L_26_0,
        F2A_L_25_6,
        F2A_L_25_4,
        F2A_L_25_2,
        F2A_L_25_0,
        F2A_L_8_6,
        F2A_L_8_4,
        F2A_L_8_2,
        F2A_L_8_0,
        F2A_L_6_15,
        F2A_L_6_13,
        F2A_L_6_11,
        F2A_L_6_9,
        F2A_L_6_6,
        F2A_L_6_4,
        F2A_L_6_2,
        F2A_L_6_0,
        F2A_L_5_9,
        F2A_L_5_7,
        F2A_L_5_5,
        F2A_L_5_3,
        F2A_L_5_0,
        F2A_L_4_13,
        F2A_L_4_11,
        F2A_L_4_9,
        F2A_L_4_6,
        F2A_L_4_4,
        F2A_L_4_2,
        F2A_L_4_0,
        F2A_L_3_6,
        F2A_L_3_4,
        F2A_L_3_2,
        F2A_L_3_0,
        F2A_L_2_6,
        F2A_L_2_4,
        F2A_L_2_2,
        F2A_L_2_0
      }),
      .lint_ADDR({
        A2F_L_15_5,
        A2F_L_15_4,
        A2F_L_15_3,
        A2F_L_15_2,
        A2F_L_15_1,
        A2F_L_15_0,
        A2F_L_14_7,
        A2F_L_14_6,
        A2F_L_14_5,
        A2F_L_14_4,
        A2F_L_14_3,
        A2F_L_14_2,
        A2F_L_14_1,
        A2F_L_14_0,
        A2F_L_13_5,
        A2F_L_13_4,
        A2F_L_13_3,
        A2F_L_13_2,
        A2F_L_13_1,
        A2F_L_13_0
      }),
      .lint_BE({A2F_L_12_7, A2F_L_12_6, A2F_L_12_5, A2F_L_12_4}),
      .lint_RDATA({
        F2A_L_15_7,
        F2A_L_15_6,
        F2A_L_15_5,
        F2A_L_15_4,
        F2A_L_15_3,
        F2A_L_15_2,
        F2A_L_15_1,
        F2A_L_15_0,
        F2A_L_14_8,
        F2A_L_14_7,
        F2A_L_14_6,
        F2A_L_14_5,
        F2A_L_14_4,
        F2A_L_14_3,
        F2A_L_14_2,
        F2A_L_14_1,
        F2A_L_13_6,
        F2A_L_13_5,
        F2A_L_13_4,
        F2A_L_13_3,
        F2A_L_13_2,
        F2A_L_13_1,
        F2A_L_13_0,
        F2A_L_12_16,
        F2A_L_12_15,
        F2A_L_12_14,
        F2A_L_12_13,
        F2A_L_12_12,
        F2A_L_12_11,
        F2A_L_12_10,
        F2A_L_12_9,
        F2A_L_12_8
      }),
      .lint_WDATA({
        A2F_L_12_1,
        A2F_L_12_0,
        A2F_L_11_5,
        A2F_L_11_4,
        A2F_L_11_3,
        A2F_L_11_2,
        A2F_L_11_1,
        A2F_L_11_0,
        A2F_L_10_7,
        A2F_L_10_6,
        A2F_L_10_5,
        A2F_L_10_4,
        A2F_L_10_3,
        A2F_L_10_2,
        A2F_L_10_1,
        A2F_L_10_0,
        A2F_L_9_5,
        A2F_L_9_4,
        A2F_L_9_3,
        A2F_L_9_2,
        A2F_L_9_1,
        A2F_L_9_0,
        A2F_L_8_7,
        A2F_L_8_6,
        A2F_L_8_5,
        A2F_L_8_4,
        A2F_L_8_3,
        A2F_L_8_2,
        A2F_L_8_1,
        A2F_L_8_0,
        A2F_L_7_5,
        A2F_L_7_4
      }),
      .m0_coef_raddr({
        F2A_T_14_14,
        F2A_T_14_15,
        F2A_T_14_16,
        F2A_T_14_17,
        F2A_T_15_1,
        F2A_T_15_2,
        F2A_T_15_3,
        F2A_T_15_4,
        F2A_T_15_5,
        F2A_T_15_6,
        F2A_T_15_7,
        F2A_T_15_8
      }),
      .m0_coef_rdata({
        A2F_T_11_4,
        A2F_T_11_5,
        A2F_T_12_0,
        A2F_T_12_1,
        A2F_T_12_2,
        A2F_T_12_3,
        A2F_T_12_4,
        A2F_T_12_5,
        A2F_T_12_6,
        A2F_T_12_7,
        A2F_T_13_0,
        A2F_T_13_1,
        A2F_T_13_2,
        A2F_T_13_3,
        A2F_T_13_4,
        A2F_T_13_5,
        A2F_T_14_0,
        A2F_T_14_1,
        A2F_T_14_2,
        A2F_T_14_3,
        A2F_T_14_4,
        A2F_T_14_5,
        A2F_T_14_6,
        A2F_T_14_7,
        A2F_T_15_0,
        A2F_T_15_1,
        A2F_T_15_2,
        A2F_T_15_3,
        A2F_T_15_4,
        A2F_T_15_5,
        A2F_T_16_0,
        A2F_T_16_1
      }),
      .m0_coef_rmode({F2A_T_14_12, F2A_T_14_13}),
      .m0_coef_waddr({
        F2A_T_13_10,
        F2A_T_13_11,
        F2A_T_14_0,
        F2A_T_14_1,
        F2A_T_14_2,
        F2A_T_14_3,
        F2A_T_14_4,
        F2A_T_14_5,
        F2A_T_14_6,
        F2A_T_14_7,
        F2A_T_14_8,
        F2A_T_14_9
      }),
      .m0_coef_wdata({
        F2A_T_11_7,
        F2A_T_11_8,
        F2A_T_11_9,
        F2A_T_11_10,
        F2A_T_11_11,
        F2A_T_12_0,
        F2A_T_12_1,
        F2A_T_12_2,
        F2A_T_12_3,
        F2A_T_12_4,
        F2A_T_12_5,
        F2A_T_12_6,
        F2A_T_12_7,
        F2A_T_12_8,
        F2A_T_12_9,
        F2A_T_12_10,
        F2A_T_12_11,
        F2A_T_12_12,
        F2A_T_12_13,
        F2A_T_12_14,
        F2A_T_12_15,
        F2A_T_12_16,
        F2A_T_12_17,
        F2A_T_13_1,
        F2A_T_13_2,
        F2A_T_13_3,
        F2A_T_13_4,
        F2A_T_13_5,
        F2A_T_13_6,
        F2A_T_13_7,
        F2A_T_13_8,
        F2A_T_13_9
      }),
      .m0_coef_wmode({F2A_T_15_9, F2A_T_15_10}),
      .m0_m0_coef_in({
        F2A_T_9_1,
        F2A_T_9_2,
        F2A_T_9_3,
        F2A_T_9_4,
        F2A_T_9_5,
        F2A_T_9_6,
        F2A_T_9_7,
        F2A_T_9_8,
        F2A_T_9_9,
        F2A_T_9_10,
        F2A_T_9_11,
        F2A_T_10_0,
        F2A_T_10_1,
        F2A_T_10_2,
        F2A_T_10_3,
        F2A_T_10_4,
        F2A_T_10_5,
        F2A_T_10_6,
        F2A_T_10_7,
        F2A_T_10_8,
        F2A_T_10_9,
        F2A_T_10_10,
        F2A_T_10_11,
        F2A_T_10_12,
        F2A_T_10_13,
        F2A_T_10_14,
        F2A_T_10_15,
        F2A_T_10_16,
        F2A_T_10_17,
        F2A_T_11_0,
        F2A_T_11_1,
        F2A_T_11_2
      }),
      .m0_m0_dataout({
        A2F_T_7_0,
        A2F_T_7_1,
        A2F_T_7_2,
        A2F_T_7_3,
        A2F_T_7_4,
        A2F_T_7_5,
        A2F_T_8_0,
        A2F_T_8_1,
        A2F_T_8_2,
        A2F_T_8_3,
        A2F_T_8_4,
        A2F_T_8_5,
        A2F_T_8_6,
        A2F_T_8_7,
        A2F_T_9_0,
        A2F_T_9_1,
        A2F_T_9_2,
        A2F_T_9_3,
        A2F_T_9_4,
        A2F_T_9_5,
        A2F_T_10_0,
        A2F_T_10_1,
        A2F_T_10_2,
        A2F_T_10_3,
        A2F_T_10_4,
        A2F_T_10_5,
        A2F_T_10_6,
        A2F_T_10_7,
        A2F_T_11_0,
        A2F_T_11_1,
        A2F_T_11_2,
        A2F_T_11_3
      }),
      .m0_m0_mode({F2A_T_11_3, F2A_T_11_4}),
      .m0_m0_oper_in({
        F2A_T_6_15,
        F2A_T_6_16,
        F2A_T_6_17,
        F2A_T_7_1,
        F2A_T_7_2,
        F2A_T_7_3,
        F2A_T_7_4,
        F2A_T_7_5,
        F2A_T_7_6,
        F2A_T_7_7,
        F2A_T_7_8,
        F2A_T_7_9,
        F2A_T_7_10,
        F2A_T_7_11,
        F2A_T_8_0,
        F2A_T_8_1,
        F2A_T_8_2,
        F2A_T_8_3,
        F2A_T_8_4,
        F2A_T_8_5,
        F2A_T_8_6,
        F2A_T_8_7,
        F2A_T_8_8,
        F2A_T_8_9,
        F2A_T_8_10,
        F2A_T_8_11,
        F2A_T_8_12,
        F2A_T_8_13,
        F2A_T_8_14,
        F2A_T_8_15,
        F2A_T_8_16,
        F2A_T_8_17
      }),
      .m0_m0_outsel({F2A_T_6_6, F2A_T_6_7, F2A_T_6_8, F2A_T_6_9, F2A_T_6_10, F2A_T_6_11}),
      .m0_m1_coef_in({
        F2A_T_19_4,
        F2A_T_19_5,
        F2A_T_19_6,
        F2A_T_19_7,
        F2A_T_19_8,
        F2A_T_19_9,
        F2A_T_19_10,
        F2A_T_19_11,
        F2A_T_20_0,
        F2A_T_20_1,
        F2A_T_20_2,
        F2A_T_20_3,
        F2A_T_20_4,
        F2A_T_20_5,
        F2A_T_20_6,
        F2A_T_20_7,
        F2A_T_20_8,
        F2A_T_20_9,
        F2A_T_20_10,
        F2A_T_20_11,
        F2A_T_20_12,
        F2A_T_20_13,
        F2A_T_20_14,
        F2A_T_20_15,
        F2A_T_20_16,
        F2A_T_20_17,
        F2A_T_21_0,
        F2A_T_21_1,
        F2A_T_21_2,
        F2A_T_21_3,
        F2A_T_21_4,
        F2A_T_21_5
      }),
      .m0_m1_dataout({
        A2F_T_18_0,
        A2F_T_18_1,
        A2F_T_18_2,
        A2F_T_18_3,
        A2F_T_18_4,
        A2F_T_18_5,
        A2F_T_18_6,
        A2F_T_18_7,
        A2F_T_19_0,
        A2F_T_19_1,
        A2F_T_19_2,
        A2F_T_19_3,
        A2F_T_19_4,
        A2F_T_19_5,
        A2F_T_20_0,
        A2F_T_20_1,
        A2F_T_20_2,
        A2F_T_20_3,
        A2F_T_20_4,
        A2F_T_20_5,
        A2F_T_20_6,
        A2F_T_21_0,
        A2F_T_21_1,
        A2F_T_21_2,
        A2F_T_21_3,
        A2F_T_21_4,
        A2F_T_21_5,
        A2F_T_22_0,
        A2F_T_22_1,
        A2F_T_22_2,
        A2F_T_22_3,
        A2F_T_22_4
      }),
      .m0_m1_mode({F2A_T_21_6, F2A_T_21_8}),
      .m0_m1_oper_in({
        F2A_T_21_9,
        F2A_T_21_10,
        F2A_T_21_11,
        F2A_T_22_0,
        F2A_T_22_1,
        F2A_T_22_2,
        F2A_T_22_3,
        F2A_T_22_4,
        F2A_T_22_5,
        F2A_T_22_6,
        F2A_T_22_7,
        F2A_T_22_8,
        F2A_T_22_9,
        F2A_T_22_10,
        F2A_T_22_11,
        F2A_T_22_12,
        F2A_T_22_13,
        F2A_T_22_14,
        F2A_T_22_15,
        F2A_T_22_16,
        F2A_T_22_17,
        F2A_T_23_0,
        F2A_T_23_1,
        F2A_T_23_2,
        F2A_T_23_3,
        F2A_T_23_4,
        F2A_T_23_5,
        F2A_T_23_6,
        F2A_T_23_7,
        F2A_T_23_8,
        F2A_T_23_9,
        F2A_T_23_10
      }),
      .m0_m1_outsel({F2A_T_18_8, F2A_T_18_9, F2A_T_18_10, F2A_T_18_11, F2A_T_18_12, F2A_T_18_13}),
      .m0_oper0_raddr({
        F2A_T_5_3,
        F2A_T_5_4,
        F2A_T_5_5,
        F2A_T_5_6,
        F2A_T_5_7,
        F2A_T_5_8,
        F2A_T_5_9,
        F2A_T_5_10,
        F2A_T_5_11,
        F2A_T_6_1,
        F2A_T_6_2,
        F2A_T_6_3
      }),
      .m0_oper0_rdata({
        A2F_T_2_0,
        A2F_T_2_1,
        A2F_T_2_2,
        A2F_T_2_3,
        A2F_T_3_0,
        A2F_T_3_1,
        A2F_T_3_2,
        A2F_T_3_3,
        A2F_T_3_4,
        A2F_T_3_5,
        A2F_T_4_0,
        A2F_T_4_1,
        A2F_T_4_2,
        A2F_T_4_3,
        A2F_T_4_4,
        A2F_T_4_5,
        A2F_T_4_6,
        A2F_T_4_7,
        A2F_T_5_0,
        A2F_T_5_1,
        A2F_T_5_2,
        A2F_T_5_3,
        A2F_T_5_4,
        A2F_T_5_5,
        A2F_T_6_0,
        A2F_T_6_1,
        A2F_T_6_2,
        A2F_T_6_3,
        A2F_T_6_4,
        A2F_T_6_5,
        A2F_T_6_6,
        A2F_T_6_7
      }),
      .m0_oper0_rmode({F2A_T_2_4, F2A_T_2_5}),
      .m0_oper0_waddr({
        F2A_T_4_8,
        F2A_T_4_9,
        F2A_T_4_10,
        F2A_T_4_11,
        F2A_T_4_12,
        F2A_T_4_13,
        F2A_T_4_14,
        F2A_T_4_15,
        F2A_T_4_16,
        F2A_T_4_17,
        F2A_T_5_0,
        F2A_T_5_1
      }),
      .m0_oper0_wdata({
        F2A_T_2_6,
        F2A_T_2_7,
        F2A_T_2_8,
        F2A_T_2_9,
        F2A_T_2_10,
        F2A_T_2_11,
        F2A_T_2_12,
        F2A_T_2_13,
        F2A_T_2_14,
        F2A_T_2_15,
        F2A_T_2_16,
        F2A_T_2_17,
        F2A_T_3_0,
        F2A_T_3_1,
        F2A_T_3_2,
        F2A_T_3_3,
        F2A_T_3_4,
        F2A_T_3_5,
        F2A_T_3_6,
        F2A_T_3_7,
        F2A_T_3_8,
        F2A_T_3_9,
        F2A_T_3_10,
        F2A_T_3_11,
        F2A_T_4_0,
        F2A_T_4_1,
        F2A_T_4_2,
        F2A_T_4_3,
        F2A_T_4_4,
        F2A_T_4_5,
        F2A_T_4_6,
        F2A_T_4_7
      }),
      .m0_oper0_wmode({F2A_T_2_1, F2A_T_2_2}),
      .m0_oper1_raddr({
        F2A_T_28_17,
        F2A_T_29_1,
        F2A_T_29_2,
        F2A_T_29_3,
        F2A_T_29_4,
        F2A_T_29_5,
        F2A_T_29_6,
        F2A_T_29_7,
        F2A_T_29_8,
        F2A_T_29_9,
        F2A_T_29_10,
        F2A_T_29_11
      }),
      .m0_oper1_rdata({
        A2F_T_25_1,
        A2F_T_25_2,
        A2F_T_25_3,
        A2F_T_25_4,
        A2F_T_25_5,
        A2F_T_26_0,
        A2F_T_26_1,
        A2F_T_26_2,
        A2F_T_26_3,
        A2F_T_26_4,
        A2F_T_26_5,
        A2F_T_26_6,
        A2F_T_26_7,
        A2F_T_27_0,
        A2F_T_27_1,
        A2F_T_27_2,
        A2F_T_27_3,
        A2F_T_27_4,
        A2F_T_27_5,
        A2F_T_28_1,
        A2F_T_28_2,
        A2F_T_28_3,
        A2F_T_28_4,
        A2F_T_28_5,
        A2F_T_28_6,
        A2F_T_28_7,
        A2F_T_29_0,
        A2F_T_29_1,
        A2F_T_29_2,
        A2F_T_29_3,
        A2F_T_29_4,
        A2F_T_29_5
      }),
      .m0_oper1_rmode({F2A_T_28_15, F2A_T_28_16}),
      .m0_oper1_waddr({
        F2A_T_27_0,
        F2A_T_27_1,
        F2A_T_27_2,
        F2A_T_27_3,
        F2A_T_27_4,
        F2A_T_27_5,
        F2A_T_27_6,
        F2A_T_27_7,
        F2A_T_27_8,
        F2A_T_27_9,
        F2A_T_27_10,
        F2A_T_27_11
      }),
      .m0_oper1_wdata({
        F2A_T_24_16,
        F2A_T_24_17,
        F2A_T_25_0,
        F2A_T_25_1,
        F2A_T_25_2,
        F2A_T_25_3,
        F2A_T_25_4,
        F2A_T_25_5,
        F2A_T_25_6,
        F2A_T_25_7,
        F2A_T_25_8,
        F2A_T_25_9,
        F2A_T_25_10,
        F2A_T_25_11,
        F2A_T_26_0,
        F2A_T_26_1,
        F2A_T_26_2,
        F2A_T_26_3,
        F2A_T_26_4,
        F2A_T_26_5,
        F2A_T_26_6,
        F2A_T_26_7,
        F2A_T_26_8,
        F2A_T_26_9,
        F2A_T_26_10,
        F2A_T_26_11,
        F2A_T_26_12,
        F2A_T_26_13,
        F2A_T_26_14,
        F2A_T_26_15,
        F2A_T_26_16,
        F2A_T_26_17
      }),
      .m0_oper1_wmode({F2A_T_28_1, F2A_T_28_2}),
      .m1_coef_raddr({
        F2A_B_14_14,
        F2A_B_14_15,
        F2A_B_14_16,
        F2A_B_14_17,
        F2A_B_15_1,
        F2A_B_15_2,
        F2A_B_15_3,
        F2A_B_15_4,
        F2A_B_15_5,
        F2A_B_15_6,
        F2A_B_15_7,
        F2A_B_15_8
      }),
      .m1_coef_rdata({
        A2F_B_11_4,
        A2F_B_11_5,
        A2F_B_12_0,
        A2F_B_12_1,
        A2F_B_12_2,
        A2F_B_12_3,
        A2F_B_12_4,
        A2F_B_12_5,
        A2F_B_12_6,
        A2F_B_12_7,
        A2F_B_13_0,
        A2F_B_13_1,
        A2F_B_13_2,
        A2F_B_13_3,
        A2F_B_13_4,
        A2F_B_13_5,
        A2F_B_14_0,
        A2F_B_14_1,
        A2F_B_14_2,
        A2F_B_14_3,
        A2F_B_14_4,
        A2F_B_14_5,
        A2F_B_14_6,
        A2F_B_14_7,
        A2F_B_15_0,
        A2F_B_15_1,
        A2F_B_15_2,
        A2F_B_15_3,
        A2F_B_15_4,
        A2F_B_15_5,
        A2F_B_16_0,
        A2F_B_16_1
      }),
      .m1_coef_rmode({F2A_B_14_12, F2A_B_14_13}),
      .m1_coef_waddr({
        F2A_B_13_10,
        F2A_B_13_11,
        F2A_B_14_0,
        F2A_B_14_1,
        F2A_B_14_2,
        F2A_B_14_3,
        F2A_B_14_4,
        F2A_B_14_5,
        F2A_B_14_6,
        F2A_B_14_7,
        F2A_B_14_8,
        F2A_B_14_9
      }),
      .m1_coef_wdata({
        F2A_B_11_7,
        F2A_B_11_8,
        F2A_B_11_9,
        F2A_B_11_10,
        F2A_B_11_11,
        F2A_B_12_0,
        F2A_B_12_1,
        F2A_B_12_2,
        F2A_B_12_3,
        F2A_B_12_4,
        F2A_B_12_5,
        F2A_B_12_6,
        F2A_B_12_7,
        F2A_B_12_8,
        F2A_B_12_9,
        F2A_B_12_10,
        F2A_B_12_11,
        F2A_B_12_12,
        F2A_B_12_13,
        F2A_B_12_14,
        F2A_B_12_15,
        F2A_B_12_16,
        F2A_B_12_17,
        F2A_B_13_1,
        F2A_B_13_2,
        F2A_B_13_3,
        F2A_B_13_4,
        F2A_B_13_5,
        F2A_B_13_6,
        F2A_B_13_7,
        F2A_B_13_8,
        F2A_B_13_9
      }),
      .m1_coef_wmode({F2A_B_15_9, F2A_B_15_10}),
      .m1_m0_coef_in({
        F2A_B_9_1,
        F2A_B_9_2,
        F2A_B_9_3,
        F2A_B_9_4,
        F2A_B_9_5,
        F2A_B_9_6,
        F2A_B_9_7,
        F2A_B_9_8,
        F2A_B_9_9,
        F2A_B_9_10,
        F2A_B_9_11,
        F2A_B_10_0,
        F2A_B_10_1,
        F2A_B_10_2,
        F2A_B_10_3,
        F2A_B_10_4,
        F2A_B_10_5,
        F2A_B_10_6,
        F2A_B_10_7,
        F2A_B_10_8,
        F2A_B_10_9,
        F2A_B_10_10,
        F2A_B_10_11,
        F2A_B_10_12,
        F2A_B_10_13,
        F2A_B_10_14,
        F2A_B_10_15,
        F2A_B_10_16,
        F2A_B_10_17,
        F2A_B_11_0,
        F2A_B_11_1,
        F2A_B_11_2
      }),
      .m1_m0_dataout({
        A2F_B_7_0,
        A2F_B_7_1,
        A2F_B_7_2,
        A2F_B_7_3,
        A2F_B_7_4,
        A2F_B_7_5,
        A2F_B_8_0,
        A2F_B_8_1,
        A2F_B_8_2,
        A2F_B_8_3,
        A2F_B_8_4,
        A2F_B_8_5,
        A2F_B_8_6,
        A2F_B_8_7,
        A2F_B_9_0,
        A2F_B_9_1,
        A2F_B_9_2,
        A2F_B_9_3,
        A2F_B_9_4,
        A2F_B_9_5,
        A2F_B_10_0,
        A2F_B_10_1,
        A2F_B_10_2,
        A2F_B_10_3,
        A2F_B_10_4,
        A2F_B_10_5,
        A2F_B_10_6,
        A2F_B_10_7,
        A2F_B_11_0,
        A2F_B_11_1,
        A2F_B_11_2,
        A2F_B_11_3
      }),
      .m1_m0_mode({F2A_B_11_3, F2A_B_11_4}),
      .m1_m0_oper_in({
        F2A_B_6_15,
        F2A_B_6_16,
        F2A_B_6_17,
        F2A_B_7_1,
        F2A_B_7_2,
        F2A_B_7_3,
        F2A_B_7_4,
        F2A_B_7_5,
        F2A_B_7_6,
        F2A_B_7_7,
        F2A_B_7_8,
        F2A_B_7_9,
        F2A_B_7_10,
        F2A_B_7_11,
        F2A_B_8_0,
        F2A_B_8_1,
        F2A_B_8_2,
        F2A_B_8_3,
        F2A_B_8_4,
        F2A_B_8_5,
        F2A_B_8_6,
        F2A_B_8_7,
        F2A_B_8_8,
        F2A_B_8_9,
        F2A_B_8_10,
        F2A_B_8_11,
        F2A_B_8_12,
        F2A_B_8_13,
        F2A_B_8_14,
        F2A_B_8_15,
        F2A_B_8_16,
        F2A_B_8_17
      }),
      .m1_m0_outsel({F2A_B_6_6, F2A_B_6_7, F2A_B_6_8, F2A_B_6_9, F2A_B_6_10, F2A_B_6_11}),
      .m1_m1_coef_in({
        F2A_B_19_4,
        F2A_B_19_5,
        F2A_B_19_6,
        F2A_B_19_7,
        F2A_B_19_8,
        F2A_B_19_9,
        F2A_B_19_10,
        F2A_B_19_11,
        F2A_B_20_0,
        F2A_B_20_1,
        F2A_B_20_2,
        F2A_B_20_3,
        F2A_B_20_4,
        F2A_B_20_5,
        F2A_B_20_6,
        F2A_B_20_7,
        F2A_B_20_8,
        F2A_B_20_9,
        F2A_B_20_10,
        F2A_B_20_11,
        F2A_B_20_12,
        F2A_B_20_13,
        F2A_B_20_14,
        F2A_B_20_15,
        F2A_B_20_16,
        F2A_B_20_17,
        F2A_B_21_0,
        F2A_B_21_1,
        F2A_B_21_2,
        F2A_B_21_3,
        F2A_B_21_4,
        F2A_B_21_5
      }),
      .m1_m1_dataout({
        A2F_B_18_6,
        A2F_B_18_7,
        A2F_B_19_0,
        A2F_B_19_1,
        A2F_B_19_2,
        A2F_B_19_3,
        A2F_B_19_4,
        A2F_B_19_5,
        A2F_B_20_0,
        A2F_B_20_1,
        A2F_B_20_2,
        A2F_B_20_3,
        A2F_B_20_4,
        A2F_B_20_5,
        A2F_B_20_6,
        A2F_B_21_0,
        A2F_B_21_1,
        A2F_B_21_2,
        A2F_B_21_3,
        A2F_B_21_4,
        A2F_B_21_5,
        A2F_B_22_0,
        A2F_B_22_1,
        A2F_B_22_2,
        A2F_B_22_3,
        A2F_B_22_4,
        A2F_B_22_5,
        A2F_B_23_0,
        A2F_B_23_1,
        A2F_B_23_2,
        A2F_B_23_3,
        A2F_B_23_4
      }),
      .m1_m1_mode({F2A_B_21_6, F2A_B_21_8}),
      .m1_m1_oper_in({
        F2A_B_21_9,
        F2A_B_21_10,
        F2A_B_21_11,
        F2A_B_22_0,
        F2A_B_22_1,
        F2A_B_22_2,
        F2A_B_22_3,
        F2A_B_22_4,
        F2A_B_22_5,
        F2A_B_22_6,
        F2A_B_22_7,
        F2A_B_22_8,
        F2A_B_22_9,
        F2A_B_22_10,
        F2A_B_22_11,
        F2A_B_22_12,
        F2A_B_22_13,
        F2A_B_22_14,
        F2A_B_22_15,
        F2A_B_22_16,
        F2A_B_22_17,
        F2A_B_23_0,
        F2A_B_23_1,
        F2A_B_23_2,
        F2A_B_23_3,
        F2A_B_23_4,
        F2A_B_23_5,
        F2A_B_23_6,
        F2A_B_23_7,
        F2A_B_23_8,
        F2A_B_23_9,
        F2A_B_23_10
      }),
      .m1_m1_outsel({F2A_B_18_7, F2A_B_18_8, F2A_B_18_9, F2A_B_18_10, F2A_B_18_11, F2A_B_18_12}),
      .m1_oper0_raddr({
        F2A_B_5_3,
        F2A_B_5_4,
        F2A_B_5_5,
        F2A_B_5_6,
        F2A_B_5_7,
        F2A_B_5_8,
        F2A_B_5_9,
        F2A_B_5_10,
        F2A_B_5_11,
        F2A_B_6_1,
        F2A_B_6_2,
        F2A_B_6_3
      }),
      .m1_oper0_rdata({
        A2F_B_2_0,
        A2F_B_2_1,
        A2F_B_2_2,
        A2F_B_2_3,
        A2F_B_3_0,
        A2F_B_3_1,
        A2F_B_3_2,
        A2F_B_3_3,
        A2F_B_3_4,
        A2F_B_3_5,
        A2F_B_4_0,
        A2F_B_4_1,
        A2F_B_4_2,
        A2F_B_4_3,
        A2F_B_4_4,
        A2F_B_4_5,
        A2F_B_4_6,
        A2F_B_4_7,
        A2F_B_5_0,
        A2F_B_5_1,
        A2F_B_5_2,
        A2F_B_5_3,
        A2F_B_5_4,
        A2F_B_5_5,
        A2F_B_6_0,
        A2F_B_6_1,
        A2F_B_6_2,
        A2F_B_6_3,
        A2F_B_6_4,
        A2F_B_6_5,
        A2F_B_6_6,
        A2F_B_6_7
      }),
      .m1_oper0_rmode({F2A_B_2_4, F2A_B_2_5}),
      .m1_oper0_waddr({
        F2A_B_4_8,
        F2A_B_4_9,
        F2A_B_4_10,
        F2A_B_4_11,
        F2A_B_4_12,
        F2A_B_4_13,
        F2A_B_4_14,
        F2A_B_4_15,
        F2A_B_4_16,
        F2A_B_4_17,
        F2A_B_5_0,
        F2A_B_5_1
      }),
      .m1_oper0_wdata({
        F2A_B_2_6,
        F2A_B_2_7,
        F2A_B_2_8,
        F2A_B_2_9,
        F2A_B_2_10,
        F2A_B_2_11,
        F2A_B_2_12,
        F2A_B_2_13,
        F2A_B_2_14,
        F2A_B_2_15,
        F2A_B_2_16,
        F2A_B_2_17,
        F2A_B_3_0,
        F2A_B_3_1,
        F2A_B_3_2,
        F2A_B_3_3,
        F2A_B_3_4,
        F2A_B_3_5,
        F2A_B_3_6,
        F2A_B_3_7,
        F2A_B_3_8,
        F2A_B_3_9,
        F2A_B_3_10,
        F2A_B_3_11,
        F2A_B_4_0,
        F2A_B_4_1,
        F2A_B_4_2,
        F2A_B_4_3,
        F2A_B_4_4,
        F2A_B_4_5,
        F2A_B_4_6,
        F2A_B_4_7
      }),
      .m1_oper0_wmode({F2A_B_2_1, F2A_B_2_2}),
      .m1_oper1_raddr({
        F2A_B_28_17,
        F2A_B_29_1,
        F2A_B_29_2,
        F2A_B_29_3,
        F2A_B_29_4,
        F2A_B_29_5,
        F2A_B_29_6,
        F2A_B_29_7,
        F2A_B_29_8,
        F2A_B_29_9,
        F2A_B_29_10,
        F2A_B_29_11
      }),
      .m1_oper1_rdata({
        A2F_B_25_1,
        A2F_B_25_2,
        A2F_B_25_3,
        A2F_B_25_4,
        A2F_B_25_5,
        A2F_B_26_0,
        A2F_B_26_1,
        A2F_B_26_2,
        A2F_B_26_3,
        A2F_B_26_4,
        A2F_B_26_5,
        A2F_B_26_6,
        A2F_B_26_7,
        A2F_B_27_0,
        A2F_B_27_1,
        A2F_B_27_2,
        A2F_B_27_3,
        A2F_B_27_4,
        A2F_B_27_5,
        A2F_B_28_1,
        A2F_B_28_2,
        A2F_B_28_3,
        A2F_B_28_4,
        A2F_B_28_5,
        A2F_B_28_6,
        A2F_B_28_7,
        A2F_B_29_0,
        A2F_B_29_1,
        A2F_B_29_2,
        A2F_B_29_3,
        A2F_B_29_4,
        A2F_B_29_5
      }),
      .m1_oper1_rmode({F2A_B_28_15, F2A_B_28_16}),
      .m1_oper1_waddr({
        F2A_B_27_0,
        F2A_B_27_1,
        F2A_B_27_2,
        F2A_B_27_3,
        F2A_B_27_4,
        F2A_B_27_5,
        F2A_B_27_6,
        F2A_B_27_7,
        F2A_B_27_8,
        F2A_B_27_9,
        F2A_B_27_10,
        F2A_B_27_11
      }),
      .m1_oper1_wdata({
        F2A_B_24_16,
        F2A_B_24_17,
        F2A_B_25_0,
        F2A_B_25_1,
        F2A_B_25_2,
        F2A_B_25_3,
        F2A_B_25_4,
        F2A_B_25_5,
        F2A_B_25_6,
        F2A_B_25_7,
        F2A_B_25_8,
        F2A_B_25_9,
        F2A_B_25_10,
        F2A_B_25_11,
        F2A_B_26_0,
        F2A_B_26_1,
        F2A_B_26_2,
        F2A_B_26_3,
        F2A_B_26_4,
        F2A_B_26_5,
        F2A_B_26_6,
        F2A_B_26_7,
        F2A_B_26_8,
        F2A_B_26_9,
        F2A_B_26_10,
        F2A_B_26_11,
        F2A_B_26_12,
        F2A_B_26_13,
        F2A_B_26_14,
        F2A_B_26_15,
        F2A_B_26_16,
        F2A_B_26_17
      }),
      .m1_oper1_wmode({F2A_B_28_1, F2A_B_28_2}),
      .status_out({
        F2A_L_22_1,
        F2A_L_22_0,
        F2A_L_21_11,
        F2A_L_21_10,
        F2A_L_21_9,
        F2A_L_21_8,
        F2A_L_21_7,
        F2A_L_21_6,
        F2A_L_21_5,
        F2A_L_21_4,
        F2A_L_21_3,
        F2A_L_21_2,
        F2A_L_21_1,
        F2A_L_21_0,
        F2A_L_20_17,
        F2A_L_20_16,
        F2A_L_20_15,
        F2A_L_20_14,
        F2A_L_20_13,
        F2A_L_20_12,
        F2A_L_20_11,
        F2A_L_20_10,
        F2A_L_20_9,
        F2A_L_20_8,
        F2A_L_20_7,
        F2A_L_20_6,
        F2A_L_20_5,
        F2A_L_20_4,
        F2A_L_20_3,
        F2A_L_20_2,
        F2A_L_20_1,
        F2A_L_20_0
      }),
      .tcdm_addr_p0({
        F2A_R_6_17,
        F2A_R_6_16,
        F2A_R_6_15,
        F2A_R_6_14,
        F2A_R_6_13,
        F2A_R_6_12,
        F2A_R_5_11,
        F2A_R_5_10,
        F2A_R_5_9,
        F2A_R_5_8,
        F2A_R_4_14,
        F2A_R_4_13,
        F2A_R_4_12,
        F2A_R_4_11,
        F2A_R_4_10,
        F2A_R_4_9,
        F2A_R_3_11,
        F2A_R_3_10,
        F2A_R_3_9,
        F2A_R_3_8
      }),
      .tcdm_addr_p1({
        F2A_R_12_17,
        F2A_R_12_16,
        F2A_R_12_15,
        F2A_R_12_14,
        F2A_R_12_13,
        F2A_R_12_12,
        F2A_R_11_11,
        F2A_R_11_10,
        F2A_R_11_9,
        F2A_R_11_8,
        F2A_R_10_14,
        F2A_R_10_13,
        F2A_R_10_12,
        F2A_R_10_11,
        F2A_R_10_10,
        F2A_R_10_9,
        F2A_R_9_11,
        F2A_R_9_10,
        F2A_R_9_9,
        F2A_R_9_8
      }),
      .tcdm_addr_p2({
        F2A_R_20_17,
        F2A_R_20_16,
        F2A_R_20_15,
        F2A_R_20_14,
        F2A_R_20_13,
        F2A_R_20_12,
        F2A_R_19_11,
        F2A_R_19_10,
        F2A_R_19_9,
        F2A_R_19_8,
        F2A_R_18_14,
        F2A_R_18_13,
        F2A_R_18_12,
        F2A_R_18_11,
        F2A_R_18_10,
        F2A_R_18_9,
        F2A_R_17_11,
        F2A_R_17_10,
        F2A_R_17_9,
        F2A_R_17_8
      }),
      .tcdm_addr_p3({
        F2A_R_26_17,
        F2A_R_26_16,
        F2A_R_26_15,
        F2A_R_26_14,
        F2A_R_26_13,
        F2A_R_26_12,
        F2A_R_25_11,
        F2A_R_25_10,
        F2A_R_25_9,
        F2A_R_25_8,
        F2A_R_24_14,
        F2A_R_24_13,
        F2A_R_24_12,
        F2A_R_24_11,
        F2A_R_24_10,
        F2A_R_24_9,
        F2A_R_23_11,
        F2A_R_23_10,
        F2A_R_23_9,
        F2A_R_23_8
      }),
      .tcdm_be_p0({F2A_R_3_6, F2A_R_3_5, F2A_R_3_4, F2A_R_3_3}),
      .tcdm_be_p1({F2A_R_9_6, F2A_R_9_5, F2A_R_9_4, F2A_R_9_3}),
      .tcdm_be_p2({F2A_R_17_6, F2A_R_17_5, F2A_R_17_4, F2A_R_17_3}),
      .tcdm_be_p3({F2A_R_23_6, F2A_R_23_5, F2A_R_23_4, F2A_R_23_3}),
      .tcdm_rdata_p0({
        A2F_R_8_3,
        A2F_R_8_2,
        A2F_R_8_1,
        A2F_R_8_0,
        A2F_R_7_5,
        A2F_R_7_4,
        A2F_R_7_3,
        A2F_R_7_2,
        A2F_R_7_1,
        A2F_R_7_0,
        A2F_R_6_6,
        A2F_R_6_5,
        A2F_R_6_4,
        A2F_R_6_3,
        A2F_R_6_2,
        A2F_R_6_1,
        A2F_R_5_3,
        A2F_R_5_2,
        A2F_R_5_1,
        A2F_R_5_0,
        A2F_R_4_7,
        A2F_R_4_6,
        A2F_R_4_5,
        A2F_R_4_4,
        A2F_R_4_3,
        A2F_R_4_2,
        A2F_R_4_1,
        A2F_R_4_0,
        A2F_R_3_3,
        A2F_R_3_2,
        A2F_R_3_1,
        A2F_R_3_0
      }),
      .tcdm_rdata_p1({
        A2F_R_14_3,
        A2F_R_14_2,
        A2F_R_14_1,
        A2F_R_14_0,
        A2F_R_13_5,
        A2F_R_13_4,
        A2F_R_13_3,
        A2F_R_13_2,
        A2F_R_13_1,
        A2F_R_13_0,
        A2F_R_12_6,
        A2F_R_12_5,
        A2F_R_12_4,
        A2F_R_12_3,
        A2F_R_12_2,
        A2F_R_12_1,
        A2F_R_11_3,
        A2F_R_11_2,
        A2F_R_11_1,
        A2F_R_11_0,
        A2F_R_10_7,
        A2F_R_10_6,
        A2F_R_10_5,
        A2F_R_10_4,
        A2F_R_10_3,
        A2F_R_10_2,
        A2F_R_10_1,
        A2F_R_10_0,
        A2F_R_9_3,
        A2F_R_9_2,
        A2F_R_9_1,
        A2F_R_9_0
      }),
      .tcdm_rdata_p2({
        A2F_R_22_3,
        A2F_R_22_2,
        A2F_R_22_1,
        A2F_R_22_0,
        A2F_R_21_5,
        A2F_R_21_4,
        A2F_R_21_3,
        A2F_R_21_2,
        A2F_R_21_1,
        A2F_R_21_0,
        A2F_R_20_6,
        A2F_R_20_5,
        A2F_R_20_4,
        A2F_R_20_3,
        A2F_R_20_2,
        A2F_R_20_1,
        A2F_R_19_3,
        A2F_R_19_2,
        A2F_R_19_1,
        A2F_R_19_0,
        A2F_R_18_7,
        A2F_R_18_6,
        A2F_R_18_5,
        A2F_R_18_4,
        A2F_R_18_3,
        A2F_R_18_2,
        A2F_R_18_1,
        A2F_R_18_0,
        A2F_R_17_3,
        A2F_R_17_2,
        A2F_R_17_1,
        A2F_R_17_0
      }),
      .tcdm_rdata_p3({
        A2F_R_28_3,
        A2F_R_28_2,
        A2F_R_28_1,
        A2F_R_28_0,
        A2F_R_27_5,
        A2F_R_27_4,
        A2F_R_27_3,
        A2F_R_27_2,
        A2F_R_27_1,
        A2F_R_27_0,
        A2F_R_26_6,
        A2F_R_26_5,
        A2F_R_26_4,
        A2F_R_26_3,
        A2F_R_26_2,
        A2F_R_26_1,
        A2F_R_25_3,
        A2F_R_25_2,
        A2F_R_25_1,
        A2F_R_25_0,
        A2F_R_24_7,
        A2F_R_24_6,
        A2F_R_24_5,
        A2F_R_24_4,
        A2F_R_24_3,
        A2F_R_24_2,
        A2F_R_24_1,
        A2F_R_24_0,
        A2F_R_23_3,
        A2F_R_23_2,
        A2F_R_23_1,
        A2F_R_23_0
      }),
      .tcdm_wdata_p0({
        F2A_R_7_7,
        F2A_R_7_6,
        F2A_R_7_5,
        F2A_R_7_4,
        F2A_R_7_3,
        F2A_R_7_2,
        F2A_R_7_1,
        F2A_R_7_0,
        F2A_R_6_7,
        F2A_R_6_6,
        F2A_R_6_5,
        F2A_R_6_4,
        F2A_R_6_3,
        F2A_R_6_2,
        F2A_R_6_1,
        F2A_R_6_0,
        F2A_R_5_7,
        F2A_R_5_6,
        F2A_R_5_5,
        F2A_R_5_4,
        F2A_R_5_3,
        F2A_R_5_2,
        F2A_R_5_1,
        F2A_R_5_0,
        F2A_R_4_7,
        F2A_R_4_6,
        F2A_R_4_5,
        F2A_R_4_4,
        F2A_R_4_3,
        F2A_R_4_2,
        F2A_R_4_1,
        F2A_R_4_0
      }),
      .tcdm_wdata_p1({
        F2A_R_13_7,
        F2A_R_13_6,
        F2A_R_13_5,
        F2A_R_13_4,
        F2A_R_13_3,
        F2A_R_13_2,
        F2A_R_13_1,
        F2A_R_13_0,
        F2A_R_12_7,
        F2A_R_12_6,
        F2A_R_12_5,
        F2A_R_12_4,
        F2A_R_12_3,
        F2A_R_12_2,
        F2A_R_12_1,
        F2A_R_12_0,
        F2A_R_11_7,
        F2A_R_11_6,
        F2A_R_11_5,
        F2A_R_11_4,
        F2A_R_11_3,
        F2A_R_11_2,
        F2A_R_11_1,
        F2A_R_11_0,
        F2A_R_10_7,
        F2A_R_10_6,
        F2A_R_10_5,
        F2A_R_10_4,
        F2A_R_10_3,
        F2A_R_10_2,
        F2A_R_10_1,
        F2A_R_10_0
      }),
      .tcdm_wdata_p2({
        F2A_R_21_7,
        F2A_R_21_6,
        F2A_R_21_5,
        F2A_R_21_4,
        F2A_R_21_3,
        F2A_R_21_2,
        F2A_R_21_1,
        F2A_R_21_0,
        F2A_R_20_7,
        F2A_R_20_6,
        F2A_R_20_5,
        F2A_R_20_4,
        F2A_R_20_3,
        F2A_R_20_2,
        F2A_R_20_1,
        F2A_R_20_0,
        F2A_R_19_7,
        F2A_R_19_6,
        F2A_R_19_5,
        F2A_R_19_4,
        F2A_R_19_3,
        F2A_R_19_2,
        F2A_R_19_1,
        F2A_R_19_0,
        F2A_R_18_7,
        F2A_R_18_6,
        F2A_R_18_5,
        F2A_R_18_4,
        F2A_R_18_3,
        F2A_R_18_2,
        F2A_R_18_1,
        F2A_R_18_0
      }),
      .tcdm_wdata_p3({
        F2A_R_27_7,
        F2A_R_27_6,
        F2A_R_27_5,
        F2A_R_27_4,
        F2A_R_27_3,
        F2A_R_27_2,
        F2A_R_27_1,
        F2A_R_27_0,
        F2A_R_26_7,
        F2A_R_26_6,
        F2A_R_26_5,
        F2A_R_26_4,
        F2A_R_26_3,
        F2A_R_26_2,
        F2A_R_26_1,
        F2A_R_26_0,
        F2A_R_25_7,
        F2A_R_25_6,
        F2A_R_25_5,
        F2A_R_25_4,
        F2A_R_25_3,
        F2A_R_25_2,
        F2A_R_25_1,
        F2A_R_25_0,
        F2A_R_24_7,
        F2A_R_24_6,
        F2A_R_24_5,
        F2A_R_24_4,
        F2A_R_24_3,
        F2A_R_24_2,
        F2A_R_24_1,
        F2A_R_24_0
      }),
      .version({
        F2Adef_L_4_0,
        F2Adef_L_2_6,
        F2Adef_L_2_5,
        F2Adef_L_2_4,
        F2Adef_L_2_3,
        F2Adef_L_2_2,
        F2Adef_L_2_1,
        F2Adef_L_2_0
      })
  );


  assign BL_DOUT_0_ = 1'b0;
  assign BL_DOUT_1_ = 1'b0;
  assign BL_DOUT_2_ = 1'b0;
  assign BL_DOUT_3_ = 1'b0;
  assign BL_DOUT_4_ = 1'b0;
  assign BL_DOUT_5_ = 1'b0;
  assign BL_DOUT_6_ = 1'b0;
  assign BL_DOUT_7_ = 1'b0;
  assign BL_DOUT_8_ = 1'b0;
  assign BL_DOUT_9_ = 1'b0;
  assign BL_DOUT_10_ = 1'b0;
  assign BL_DOUT_11_ = 1'b0;
  assign BL_DOUT_12_ = 1'b0;
  assign BL_DOUT_13_ = 1'b0;
  assign BL_DOUT_14_ = 1'b0;
  assign BL_DOUT_15_ = 1'b0;
  assign BL_DOUT_16_ = 1'b0;
  assign BL_DOUT_17_ = 1'b0;
  assign BL_DOUT_18_ = 1'b0;
  assign BL_DOUT_19_ = 1'b0;
  assign BL_DOUT_20_ = 1'b0;
  assign BL_DOUT_21_ = 1'b0;
  assign BL_DOUT_22_ = 1'b0;
  assign BL_DOUT_23_ = 1'b0;
  assign BL_DOUT_24_ = 1'b0;
  assign BL_DOUT_25_ = 1'b0;
  assign BL_DOUT_26_ = 1'b0;
  assign BL_DOUT_27_ = 1'b0;
  assign BL_DOUT_28_ = 1'b0;
  assign BL_DOUT_29_ = 1'b0;
  assign BL_DOUT_30_ = 1'b0;
  assign BL_DOUT_31_ = 1'b0;
  assign FB_SPE_OUT_0_ = 1'b0;
  assign FB_SPE_OUT_1_ = 1'b0;
  assign FB_SPE_OUT_2_ = 1'b0;
  assign FB_SPE_OUT_3_ = 1'b0;
  assign PARALLEL_CFG = 1'b0;
  assign F2A_B_15_11 = 1'b0;
  assign F2A_B_16_0 = 1'b0;
  assign F2A_B_16_1 = 1'b0;
  assign F2A_B_16_10 = 1'b0;
  assign F2A_B_16_11 = 1'b0;
  assign F2A_B_16_12 = 1'b0;
  assign F2A_B_16_13 = 1'b0;
  assign F2A_B_16_17 = 1'b0;
  assign F2A_B_16_2 = 1'b0;
  assign F2A_B_16_3 = 1'b0;
  assign F2A_B_16_4 = 1'b0;
  assign F2A_B_16_5 = 1'b0;
  assign F2A_B_16_6 = 1'b0;
  assign F2A_B_16_7 = 1'b0;
  assign F2A_B_16_8 = 1'b0;
  assign F2A_B_16_9 = 1'b0;
  assign F2A_B_17_0 = 1'b0;
  assign F2A_B_17_1 = 1'b0;
  assign F2A_B_17_10 = 1'b0;
  assign F2A_B_17_11 = 1'b0;
  assign F2A_B_17_2 = 1'b0;
  assign F2A_B_17_3 = 1'b0;
  assign F2A_B_17_4 = 1'b0;
  assign F2A_B_17_5 = 1'b0;
  assign F2A_B_17_6 = 1'b0;
  assign F2A_B_17_7 = 1'b0;
  assign F2A_B_17_8 = 1'b0;
  assign F2A_B_17_9 = 1'b0;
  assign F2A_B_18_0 = 1'b0;
  assign F2A_B_18_1 = 1'b0;
  assign F2A_B_18_17 = 1'b0;
  assign F2A_B_18_2 = 1'b0;
  assign F2A_B_18_3 = 1'b0;
  assign F2A_B_18_4 = 1'b0;
  assign F2A_B_18_5 = 1'b0;
  assign F2A_B_18_6 = 1'b0;
  assign F2A_B_1_0 = 1'b0;
  assign F2A_B_1_1 = 1'b0;
  assign F2A_B_1_10 = 1'b0;
  assign F2A_B_1_11 = 1'b0;
  assign F2A_B_1_2 = 1'b0;
  assign F2A_B_1_3 = 1'b0;
  assign F2A_B_1_4 = 1'b0;
  assign F2A_B_1_5 = 1'b0;
  assign F2A_B_1_6 = 1'b0;
  assign F2A_B_1_7 = 1'b0;
  assign F2A_B_1_8 = 1'b0;
  assign F2A_B_1_9 = 1'b0;
  assign F2A_B_23_11 = 1'b0;
  assign F2A_B_24_0 = 1'b0;
  assign F2A_B_24_1 = 1'b0;
  assign F2A_B_24_10 = 1'b0;
  assign F2A_B_24_11 = 1'b0;
  assign F2A_B_24_12 = 1'b0;
  assign F2A_B_24_13 = 1'b0;
  assign F2A_B_24_14 = 1'b0;
  assign F2A_B_24_15 = 1'b0;
  assign F2A_B_24_2 = 1'b0;
  assign F2A_B_24_3 = 1'b0;
  assign F2A_B_24_4 = 1'b0;
  assign F2A_B_24_5 = 1'b0;
  assign F2A_B_24_6 = 1'b0;
  assign F2A_B_24_7 = 1'b0;
  assign F2A_B_24_8 = 1'b0;
  assign F2A_B_24_9 = 1'b0;
  assign F2A_B_28_10 = 1'b0;
  assign F2A_B_28_11 = 1'b0;
  assign F2A_B_28_12 = 1'b0;
  assign F2A_B_28_13 = 1'b0;
  assign F2A_B_28_14 = 1'b0;
  assign F2A_B_28_5 = 1'b0;
  assign F2A_B_28_6 = 1'b0;
  assign F2A_B_28_7 = 1'b0;
  assign F2A_B_28_8 = 1'b0;
  assign F2A_B_28_9 = 1'b0;
  assign F2A_B_30_0 = 1'b0;
  assign F2A_B_30_1 = 1'b0;
  assign F2A_B_30_10 = 1'b0;
  assign F2A_B_30_11 = 1'b0;
  assign F2A_B_30_12 = 1'b0;
  assign F2A_B_30_13 = 1'b0;
  assign F2A_B_30_14 = 1'b0;
  assign F2A_B_30_15 = 1'b0;
  assign F2A_B_30_16 = 1'b0;
  assign F2A_B_30_17 = 1'b0;
  assign F2A_B_30_2 = 1'b0;
  assign F2A_B_30_3 = 1'b0;
  assign F2A_B_30_4 = 1'b0;
  assign F2A_B_30_5 = 1'b0;
  assign F2A_B_30_6 = 1'b0;
  assign F2A_B_30_7 = 1'b0;
  assign F2A_B_30_8 = 1'b0;
  assign F2A_B_30_9 = 1'b0;
  assign F2A_B_31_0 = 1'b0;
  assign F2A_B_31_1 = 1'b0;
  assign F2A_B_31_10 = 1'b0;
  assign F2A_B_31_11 = 1'b0;
  assign F2A_B_31_2 = 1'b0;
  assign F2A_B_31_3 = 1'b0;
  assign F2A_B_31_4 = 1'b0;
  assign F2A_B_31_5 = 1'b0;
  assign F2A_B_31_6 = 1'b0;
  assign F2A_B_31_7 = 1'b0;
  assign F2A_B_31_8 = 1'b0;
  assign F2A_B_31_9 = 1'b0;
  assign F2A_B_32_0 = 1'b0;
  assign F2A_B_32_1 = 1'b0;
  assign F2A_B_32_10 = 1'b0;
  assign F2A_B_32_11 = 1'b0;
  assign F2A_B_32_12 = 1'b0;
  assign F2A_B_32_13 = 1'b0;
  assign F2A_B_32_14 = 1'b0;
  assign F2A_B_32_15 = 1'b0;
  assign F2A_B_32_16 = 1'b0;
  assign F2A_B_32_17 = 1'b0;
  assign F2A_B_32_2 = 1'b0;
  assign F2A_B_32_3 = 1'b0;
  assign F2A_B_32_4 = 1'b0;
  assign F2A_B_32_5 = 1'b0;
  assign F2A_B_32_6 = 1'b0;
  assign F2A_B_32_7 = 1'b0;
  assign F2A_B_32_8 = 1'b0;
  assign F2A_B_32_9 = 1'b0;
  assign F2A_L_10_0 = 1'b0;
  assign F2A_L_10_1 = 1'b0;
  assign F2A_L_10_10 = 1'b0;
  assign F2A_L_10_11 = 1'b0;
  assign F2A_L_10_12 = 1'b0;
  assign F2A_L_10_13 = 1'b0;
  assign F2A_L_10_14 = 1'b0;
  assign F2A_L_10_15 = 1'b0;
  assign F2A_L_10_16 = 1'b0;
  assign F2A_L_10_17 = 1'b0;
  assign F2A_L_10_2 = 1'b0;
  assign F2A_L_10_3 = 1'b0;
  assign F2A_L_10_4 = 1'b0;
  assign F2A_L_10_5 = 1'b0;
  assign F2A_L_10_6 = 1'b0;
  assign F2A_L_10_7 = 1'b0;
  assign F2A_L_10_8 = 1'b0;
  assign F2A_L_10_9 = 1'b0;
  assign F2A_L_11_0 = 1'b0;
  assign F2A_L_11_1 = 1'b0;
  assign F2A_L_11_10 = 1'b0;
  assign F2A_L_11_11 = 1'b0;
  assign F2A_L_11_2 = 1'b0;
  assign F2A_L_11_3 = 1'b0;
  assign F2A_L_11_4 = 1'b0;
  assign F2A_L_11_5 = 1'b0;
  assign F2A_L_11_6 = 1'b0;
  assign F2A_L_11_7 = 1'b0;
  assign F2A_L_11_8 = 1'b0;
  assign F2A_L_11_9 = 1'b0;
  assign F2A_L_12_0 = 1'b0;
  assign F2A_L_12_1 = 1'b0;
  assign F2A_L_12_17 = 1'b0;
  assign F2A_L_12_2 = 1'b0;
  assign F2A_L_12_3 = 1'b0;
  assign F2A_L_12_4 = 1'b0;
  assign F2A_L_12_5 = 1'b0;
  assign F2A_L_12_6 = 1'b0;
  assign F2A_L_12_7 = 1'b0;
  assign F2A_L_13_10 = 1'b0;
  assign F2A_L_13_11 = 1'b0;
  assign F2A_L_13_7 = 1'b0;
  assign F2A_L_13_8 = 1'b0;
  assign F2A_L_13_9 = 1'b0;
  assign F2A_L_14_10 = 1'b0;
  assign F2A_L_14_11 = 1'b0;
  assign F2A_L_14_12 = 1'b0;
  assign F2A_L_14_13 = 1'b0;
  assign F2A_L_14_14 = 1'b0;
  assign F2A_L_14_15 = 1'b0;
  assign F2A_L_14_16 = 1'b0;
  assign F2A_L_14_17 = 1'b0;
  assign F2A_L_15_10 = 1'b0;
  assign F2A_L_15_11 = 1'b0;
  assign F2A_L_15_9 = 1'b0;
  assign F2A_L_16_0 = 1'b0;
  assign F2A_L_16_1 = 1'b0;
  assign F2A_L_16_10 = 1'b0;
  assign F2A_L_16_11 = 1'b0;
  assign F2A_L_16_12 = 1'b0;
  assign F2A_L_16_13 = 1'b0;
  assign F2A_L_16_14 = 1'b0;
  assign F2A_L_16_15 = 1'b0;
  assign F2A_L_16_16 = 1'b0;
  assign F2A_L_16_17 = 1'b0;
  assign F2A_L_16_2 = 1'b0;
  assign F2A_L_16_3 = 1'b0;
  assign F2A_L_16_4 = 1'b0;
  assign F2A_L_16_5 = 1'b0;
  assign F2A_L_16_6 = 1'b0;
  assign F2A_L_16_7 = 1'b0;
  assign F2A_L_16_8 = 1'b0;
  assign F2A_L_16_9 = 1'b0;
  assign F2A_L_17_10 = 1'b0;
  assign F2A_L_17_11 = 1'b0;
  assign F2A_L_17_8 = 1'b0;
  assign F2A_L_17_9 = 1'b0;
  assign F2A_L_18_16 = 1'b0;
  assign F2A_L_18_17 = 1'b0;
  assign F2A_L_19_10 = 1'b0;
  assign F2A_L_19_11 = 1'b0;
  assign F2A_L_19_8 = 1'b0;
  assign F2A_L_19_9 = 1'b0;
  assign F2A_L_1_0 = 1'b0;
  assign F2A_L_1_1 = 1'b0;
  assign F2A_L_1_10 = 1'b0;
  assign F2A_L_1_11 = 1'b0;
  assign F2A_L_1_2 = 1'b0;
  assign F2A_L_1_3 = 1'b0;
  assign F2A_L_1_4 = 1'b0;
  assign F2A_L_1_5 = 1'b0;
  assign F2A_L_1_6 = 1'b0;
  assign F2A_L_1_7 = 1'b0;
  assign F2A_L_1_8 = 1'b0;
  assign F2A_L_1_9 = 1'b0;
  assign F2A_L_22_10 = 1'b0;
  assign F2A_L_22_11 = 1'b0;
  assign F2A_L_22_12 = 1'b0;
  assign F2A_L_22_13 = 1'b0;
  assign F2A_L_22_14 = 1'b0;
  assign F2A_L_22_15 = 1'b0;
  assign F2A_L_22_16 = 1'b0;
  assign F2A_L_22_17 = 1'b0;
  assign F2A_L_22_2 = 1'b0;
  assign F2A_L_22_3 = 1'b0;
  assign F2A_L_22_4 = 1'b0;
  assign F2A_L_22_5 = 1'b0;
  assign F2A_L_22_6 = 1'b0;
  assign F2A_L_22_7 = 1'b0;
  assign F2A_L_22_8 = 1'b0;
  assign F2A_L_22_9 = 1'b0;
  assign F2A_L_23_0 = 1'b0;
  assign F2A_L_23_1 = 1'b0;
  assign F2A_L_23_10 = 1'b0;
  assign F2A_L_23_11 = 1'b0;
  assign F2A_L_23_2 = 1'b0;
  assign F2A_L_23_3 = 1'b0;
  assign F2A_L_23_4 = 1'b0;
  assign F2A_L_23_5 = 1'b0;
  assign F2A_L_23_6 = 1'b0;
  assign F2A_L_23_7 = 1'b0;
  assign F2A_L_23_8 = 1'b0;
  assign F2A_L_23_9 = 1'b0;
  assign F2A_L_24_0 = 1'b0;
  assign F2A_L_24_1 = 1'b0;
  assign F2A_L_24_10 = 1'b0;
  assign F2A_L_24_11 = 1'b0;
  assign F2A_L_24_12 = 1'b0;
  assign F2A_L_24_13 = 1'b0;
  assign F2A_L_24_14 = 1'b0;
  assign F2A_L_24_15 = 1'b0;
  assign F2A_L_24_16 = 1'b0;
  assign F2A_L_24_17 = 1'b0;
  assign F2A_L_24_2 = 1'b0;
  assign F2A_L_24_3 = 1'b0;
  assign F2A_L_24_4 = 1'b0;
  assign F2A_L_24_5 = 1'b0;
  assign F2A_L_24_6 = 1'b0;
  assign F2A_L_24_7 = 1'b0;
  assign F2A_L_24_8 = 1'b0;
  assign F2A_L_24_9 = 1'b0;
  assign F2A_L_25_10 = 1'b0;
  assign F2A_L_25_11 = 1'b0;
  assign F2A_L_25_9 = 1'b0;
  assign F2A_L_26_10 = 1'b0;
  assign F2A_L_26_11 = 1'b0;
  assign F2A_L_26_12 = 1'b0;
  assign F2A_L_26_13 = 1'b0;
  assign F2A_L_26_14 = 1'b0;
  assign F2A_L_26_15 = 1'b0;
  assign F2A_L_26_16 = 1'b0;
  assign F2A_L_26_17 = 1'b0;
  assign F2A_L_26_9 = 1'b0;
  assign F2A_L_27_10 = 1'b0;
  assign F2A_L_27_11 = 1'b0;
  assign F2A_L_27_9 = 1'b0;
  assign F2A_L_28_10 = 1'b0;
  assign F2A_L_28_11 = 1'b0;
  assign F2A_L_28_12 = 1'b0;
  assign F2A_L_28_13 = 1'b0;
  assign F2A_L_28_14 = 1'b0;
  assign F2A_L_28_15 = 1'b0;
  assign F2A_L_28_16 = 1'b0;
  assign F2A_L_28_17 = 1'b0;
  assign F2A_L_28_9 = 1'b0;
  assign F2A_L_29_10 = 1'b0;
  assign F2A_L_29_11 = 1'b0;
  assign F2A_L_29_9 = 1'b0;
  assign F2A_L_2_10 = 1'b0;
  assign F2A_L_2_11 = 1'b0;
  assign F2A_L_2_12 = 1'b0;
  assign F2A_L_2_13 = 1'b0;
  assign F2A_L_2_14 = 1'b0;
  assign F2A_L_2_15 = 1'b0;
  assign F2A_L_2_16 = 1'b0;
  assign F2A_L_2_17 = 1'b0;
  assign F2A_L_2_9 = 1'b0;
  assign F2A_L_30_10 = 1'b0;
  assign F2A_L_30_11 = 1'b0;
  assign F2A_L_30_12 = 1'b0;
  assign F2A_L_30_13 = 1'b0;
  assign F2A_L_30_14 = 1'b0;
  assign F2A_L_30_15 = 1'b0;
  assign F2A_L_30_16 = 1'b0;
  assign F2A_L_30_17 = 1'b0;
  assign F2A_L_30_9 = 1'b0;
  assign F2A_L_31_10 = 1'b0;
  assign F2A_L_31_11 = 1'b0;
  assign F2A_L_31_9 = 1'b0;
  assign F2A_L_32_10 = 1'b0;
  assign F2A_L_32_11 = 1'b0;
  assign F2A_L_32_12 = 1'b0;
  assign F2A_L_32_13 = 1'b0;
  assign F2A_L_32_14 = 1'b0;
  assign F2A_L_32_15 = 1'b0;
  assign F2A_L_32_16 = 1'b0;
  assign F2A_L_32_17 = 1'b0;
  assign F2A_L_32_9 = 1'b0;
  assign F2A_L_3_10 = 1'b0;
  assign F2A_L_3_11 = 1'b0;
  assign F2A_L_3_9 = 1'b0;
  assign F2A_L_4_15 = 1'b0;
  assign F2A_L_4_16 = 1'b0;
  assign F2A_L_4_17 = 1'b0;
  assign F2A_L_7_0 = 1'b0;
  assign F2A_L_7_1 = 1'b0;
  assign F2A_L_7_10 = 1'b0;
  assign F2A_L_7_11 = 1'b0;
  assign F2A_L_7_2 = 1'b0;
  assign F2A_L_7_3 = 1'b0;
  assign F2A_L_7_4 = 1'b0;
  assign F2A_L_7_5 = 1'b0;
  assign F2A_L_7_6 = 1'b0;
  assign F2A_L_7_7 = 1'b0;
  assign F2A_L_7_8 = 1'b0;
  assign F2A_L_7_9 = 1'b0;
  assign F2A_L_8_10 = 1'b0;
  assign F2A_L_8_11 = 1'b0;
  assign F2A_L_8_12 = 1'b0;
  assign F2A_L_8_13 = 1'b0;
  assign F2A_L_8_14 = 1'b0;
  assign F2A_L_8_15 = 1'b0;
  assign F2A_L_8_16 = 1'b0;
  assign F2A_L_8_17 = 1'b0;
  assign F2A_L_8_9 = 1'b0;
  assign F2A_L_9_0 = 1'b0;
  assign F2A_L_9_1 = 1'b0;
  assign F2A_L_9_10 = 1'b0;
  assign F2A_L_9_11 = 1'b0;
  assign F2A_L_9_2 = 1'b0;
  assign F2A_L_9_3 = 1'b0;
  assign F2A_L_9_4 = 1'b0;
  assign F2A_L_9_5 = 1'b0;
  assign F2A_L_9_6 = 1'b0;
  assign F2A_L_9_7 = 1'b0;
  assign F2A_L_9_8 = 1'b0;
  assign F2A_L_9_9 = 1'b0;
  assign F2A_R_10_15 = 1'b0;
  assign F2A_R_10_16 = 1'b0;
  assign F2A_R_10_17 = 1'b0;
  assign F2A_R_10_8 = 1'b0;
  assign F2A_R_12_10 = 1'b0;
  assign F2A_R_12_11 = 1'b0;
  assign F2A_R_12_8 = 1'b0;
  assign F2A_R_12_9 = 1'b0;
  assign F2A_R_13_10 = 1'b0;
  assign F2A_R_13_11 = 1'b0;
  assign F2A_R_13_8 = 1'b0;
  assign F2A_R_13_9 = 1'b0;
  assign F2A_R_14_0 = 1'b0;
  assign F2A_R_14_1 = 1'b0;
  assign F2A_R_14_10 = 1'b0;
  assign F2A_R_14_11 = 1'b0;
  assign F2A_R_14_12 = 1'b0;
  assign F2A_R_14_13 = 1'b0;
  assign F2A_R_14_14 = 1'b0;
  assign F2A_R_14_15 = 1'b0;
  assign F2A_R_14_16 = 1'b0;
  assign F2A_R_14_17 = 1'b0;
  assign F2A_R_14_2 = 1'b0;
  assign F2A_R_14_3 = 1'b0;
  assign F2A_R_14_4 = 1'b0;
  assign F2A_R_14_5 = 1'b0;
  assign F2A_R_14_6 = 1'b0;
  assign F2A_R_14_7 = 1'b0;
  assign F2A_R_14_8 = 1'b0;
  assign F2A_R_14_9 = 1'b0;
  assign F2A_R_15_0 = 1'b0;
  assign F2A_R_15_1 = 1'b0;
  assign F2A_R_15_10 = 1'b0;
  assign F2A_R_15_11 = 1'b0;
  assign F2A_R_15_2 = 1'b0;
  assign F2A_R_15_3 = 1'b0;
  assign F2A_R_15_4 = 1'b0;
  assign F2A_R_15_5 = 1'b0;
  assign F2A_R_15_6 = 1'b0;
  assign F2A_R_15_7 = 1'b0;
  assign F2A_R_15_8 = 1'b0;
  assign F2A_R_15_9 = 1'b0;
  assign F2A_R_16_0 = 1'b0;
  assign F2A_R_16_1 = 1'b0;
  assign F2A_R_16_10 = 1'b0;
  assign F2A_R_16_11 = 1'b0;
  assign F2A_R_16_12 = 1'b0;
  assign F2A_R_16_13 = 1'b0;
  assign F2A_R_16_14 = 1'b0;
  assign F2A_R_16_15 = 1'b0;
  assign F2A_R_16_16 = 1'b0;
  assign F2A_R_16_17 = 1'b0;
  assign F2A_R_16_2 = 1'b0;
  assign F2A_R_16_3 = 1'b0;
  assign F2A_R_16_4 = 1'b0;
  assign F2A_R_16_5 = 1'b0;
  assign F2A_R_16_6 = 1'b0;
  assign F2A_R_16_7 = 1'b0;
  assign F2A_R_16_8 = 1'b0;
  assign F2A_R_16_9 = 1'b0;
  assign F2A_R_17_7 = 1'b0;
  assign F2A_R_18_15 = 1'b0;
  assign F2A_R_18_16 = 1'b0;
  assign F2A_R_18_17 = 1'b0;
  assign F2A_R_18_8 = 1'b0;
  assign F2A_R_1_0 = 1'b0;
  assign F2A_R_1_1 = 1'b0;
  assign F2A_R_1_10 = 1'b0;
  assign F2A_R_1_11 = 1'b0;
  assign F2A_R_1_2 = 1'b0;
  assign F2A_R_1_3 = 1'b0;
  assign F2A_R_1_4 = 1'b0;
  assign F2A_R_1_5 = 1'b0;
  assign F2A_R_1_6 = 1'b0;
  assign F2A_R_1_7 = 1'b0;
  assign F2A_R_1_8 = 1'b0;
  assign F2A_R_1_9 = 1'b0;
  assign F2A_R_20_10 = 1'b0;
  assign F2A_R_20_11 = 1'b0;
  assign F2A_R_20_8 = 1'b0;
  assign F2A_R_20_9 = 1'b0;
  assign F2A_R_21_10 = 1'b0;
  assign F2A_R_21_11 = 1'b0;
  assign F2A_R_21_8 = 1'b0;
  assign F2A_R_21_9 = 1'b0;
  assign F2A_R_22_0 = 1'b0;
  assign F2A_R_22_1 = 1'b0;
  assign F2A_R_22_10 = 1'b0;
  assign F2A_R_22_11 = 1'b0;
  assign F2A_R_22_12 = 1'b0;
  assign F2A_R_22_13 = 1'b0;
  assign F2A_R_22_14 = 1'b0;
  assign F2A_R_22_15 = 1'b0;
  assign F2A_R_22_16 = 1'b0;
  assign F2A_R_22_17 = 1'b0;
  assign F2A_R_22_2 = 1'b0;
  assign F2A_R_22_3 = 1'b0;
  assign F2A_R_22_4 = 1'b0;
  assign F2A_R_22_5 = 1'b0;
  assign F2A_R_22_6 = 1'b0;
  assign F2A_R_22_7 = 1'b0;
  assign F2A_R_22_8 = 1'b0;
  assign F2A_R_22_9 = 1'b0;
  assign F2A_R_23_7 = 1'b0;
  assign F2A_R_24_15 = 1'b0;
  assign F2A_R_24_16 = 1'b0;
  assign F2A_R_24_17 = 1'b0;
  assign F2A_R_24_8 = 1'b0;
  assign F2A_R_26_10 = 1'b0;
  assign F2A_R_26_11 = 1'b0;
  assign F2A_R_26_8 = 1'b0;
  assign F2A_R_26_9 = 1'b0;
  assign F2A_R_27_10 = 1'b0;
  assign F2A_R_27_11 = 1'b0;
  assign F2A_R_27_8 = 1'b0;
  assign F2A_R_27_9 = 1'b0;
  assign F2A_R_28_0 = 1'b0;
  assign F2A_R_28_1 = 1'b0;
  assign F2A_R_28_10 = 1'b0;
  assign F2A_R_28_11 = 1'b0;
  assign F2A_R_28_12 = 1'b0;
  assign F2A_R_28_13 = 1'b0;
  assign F2A_R_28_14 = 1'b0;
  assign F2A_R_28_15 = 1'b0;
  assign F2A_R_28_16 = 1'b0;
  assign F2A_R_28_17 = 1'b0;
  assign F2A_R_28_2 = 1'b0;
  assign F2A_R_28_3 = 1'b0;
  assign F2A_R_28_4 = 1'b0;
  assign F2A_R_28_5 = 1'b0;
  assign F2A_R_28_6 = 1'b0;
  assign F2A_R_28_7 = 1'b0;
  assign F2A_R_28_8 = 1'b0;
  assign F2A_R_28_9 = 1'b0;
  assign F2A_R_29_0 = 1'b0;
  assign F2A_R_29_1 = 1'b0;
  assign F2A_R_29_10 = 1'b0;
  assign F2A_R_29_11 = 1'b0;
  assign F2A_R_29_2 = 1'b0;
  assign F2A_R_29_3 = 1'b0;
  assign F2A_R_29_4 = 1'b0;
  assign F2A_R_29_5 = 1'b0;
  assign F2A_R_29_6 = 1'b0;
  assign F2A_R_29_7 = 1'b0;
  assign F2A_R_29_8 = 1'b0;
  assign F2A_R_29_9 = 1'b0;
  assign F2A_R_2_0 = 1'b0;
  assign F2A_R_2_1 = 1'b0;
  assign F2A_R_2_10 = 1'b0;
  assign F2A_R_2_11 = 1'b0;
  assign F2A_R_2_12 = 1'b0;
  assign F2A_R_2_13 = 1'b0;
  assign F2A_R_2_14 = 1'b0;
  assign F2A_R_2_15 = 1'b0;
  assign F2A_R_2_16 = 1'b0;
  assign F2A_R_2_17 = 1'b0;
  assign F2A_R_2_2 = 1'b0;
  assign F2A_R_2_3 = 1'b0;
  assign F2A_R_2_4 = 1'b0;
  assign F2A_R_2_5 = 1'b0;
  assign F2A_R_2_6 = 1'b0;
  assign F2A_R_2_7 = 1'b0;
  assign F2A_R_2_8 = 1'b0;
  assign F2A_R_2_9 = 1'b0;
  assign F2A_R_30_0 = 1'b0;
  assign F2A_R_30_1 = 1'b0;
  assign F2A_R_30_10 = 1'b0;
  assign F2A_R_30_11 = 1'b0;
  assign F2A_R_30_12 = 1'b0;
  assign F2A_R_30_13 = 1'b0;
  assign F2A_R_30_14 = 1'b0;
  assign F2A_R_30_15 = 1'b0;
  assign F2A_R_30_16 = 1'b0;
  assign F2A_R_30_17 = 1'b0;
  assign F2A_R_30_2 = 1'b0;
  assign F2A_R_30_3 = 1'b0;
  assign F2A_R_30_4 = 1'b0;
  assign F2A_R_30_5 = 1'b0;
  assign F2A_R_30_6 = 1'b0;
  assign F2A_R_30_7 = 1'b0;
  assign F2A_R_30_8 = 1'b0;
  assign F2A_R_30_9 = 1'b0;
  assign F2A_R_31_0 = 1'b0;
  assign F2A_R_31_1 = 1'b0;
  assign F2A_R_31_10 = 1'b0;
  assign F2A_R_31_11 = 1'b0;
  assign F2A_R_31_2 = 1'b0;
  assign F2A_R_31_3 = 1'b0;
  assign F2A_R_31_4 = 1'b0;
  assign F2A_R_31_5 = 1'b0;
  assign F2A_R_31_6 = 1'b0;
  assign F2A_R_31_7 = 1'b0;
  assign F2A_R_31_8 = 1'b0;
  assign F2A_R_31_9 = 1'b0;
  assign F2A_R_32_0 = 1'b0;
  assign F2A_R_32_1 = 1'b0;
  assign F2A_R_32_10 = 1'b0;
  assign F2A_R_32_11 = 1'b0;
  assign F2A_R_32_12 = 1'b0;
  assign F2A_R_32_13 = 1'b0;
  assign F2A_R_32_14 = 1'b0;
  assign F2A_R_32_15 = 1'b0;
  assign F2A_R_32_16 = 1'b0;
  assign F2A_R_32_17 = 1'b0;
  assign F2A_R_32_2 = 1'b0;
  assign F2A_R_32_3 = 1'b0;
  assign F2A_R_32_4 = 1'b0;
  assign F2A_R_32_5 = 1'b0;
  assign F2A_R_32_6 = 1'b0;
  assign F2A_R_32_7 = 1'b0;
  assign F2A_R_32_8 = 1'b0;
  assign F2A_R_32_9 = 1'b0;
  assign F2A_R_3_7 = 1'b0;
  assign F2A_R_4_15 = 1'b0;
  assign F2A_R_4_16 = 1'b0;
  assign F2A_R_4_17 = 1'b0;
  assign F2A_R_4_8 = 1'b0;
  assign F2A_R_6_10 = 1'b0;
  assign F2A_R_6_11 = 1'b0;
  assign F2A_R_6_8 = 1'b0;
  assign F2A_R_6_9 = 1'b0;
  assign F2A_R_7_10 = 1'b0;
  assign F2A_R_7_11 = 1'b0;
  assign F2A_R_7_8 = 1'b0;
  assign F2A_R_7_9 = 1'b0;
  assign F2A_R_8_0 = 1'b0;
  assign F2A_R_8_1 = 1'b0;
  assign F2A_R_8_10 = 1'b0;
  assign F2A_R_8_11 = 1'b0;
  assign F2A_R_8_12 = 1'b0;
  assign F2A_R_8_13 = 1'b0;
  assign F2A_R_8_14 = 1'b0;
  assign F2A_R_8_15 = 1'b0;
  assign F2A_R_8_16 = 1'b0;
  assign F2A_R_8_17 = 1'b0;
  assign F2A_R_8_2 = 1'b0;
  assign F2A_R_8_3 = 1'b0;
  assign F2A_R_8_4 = 1'b0;
  assign F2A_R_8_5 = 1'b0;
  assign F2A_R_8_6 = 1'b0;
  assign F2A_R_8_7 = 1'b0;
  assign F2A_R_8_8 = 1'b0;
  assign F2A_R_8_9 = 1'b0;
  assign F2A_R_9_7 = 1'b0;
  assign F2A_T_15_11 = 1'b0;
  assign F2A_T_16_0 = 1'b0;
  assign F2A_T_16_1 = 1'b0;
  assign F2A_T_16_10 = 1'b0;
  assign F2A_T_16_11 = 1'b0;
  assign F2A_T_16_12 = 1'b0;
  assign F2A_T_16_13 = 1'b0;
  assign F2A_T_16_17 = 1'b0;
  assign F2A_T_16_2 = 1'b0;
  assign F2A_T_16_3 = 1'b0;
  assign F2A_T_16_4 = 1'b0;
  assign F2A_T_16_5 = 1'b0;
  assign F2A_T_16_6 = 1'b0;
  assign F2A_T_16_7 = 1'b0;
  assign F2A_T_16_8 = 1'b0;
  assign F2A_T_16_9 = 1'b0;
  assign F2A_T_17_0 = 1'b0;
  assign F2A_T_17_1 = 1'b0;
  assign F2A_T_17_10 = 1'b0;
  assign F2A_T_17_11 = 1'b0;
  assign F2A_T_17_2 = 1'b0;
  assign F2A_T_17_3 = 1'b0;
  assign F2A_T_17_4 = 1'b0;
  assign F2A_T_17_5 = 1'b0;
  assign F2A_T_17_6 = 1'b0;
  assign F2A_T_17_7 = 1'b0;
  assign F2A_T_17_8 = 1'b0;
  assign F2A_T_17_9 = 1'b0;
  assign F2A_T_18_0 = 1'b0;
  assign F2A_T_18_1 = 1'b0;
  assign F2A_T_18_2 = 1'b0;
  assign F2A_T_18_3 = 1'b0;
  assign F2A_T_18_4 = 1'b0;
  assign F2A_T_18_5 = 1'b0;
  assign F2A_T_18_6 = 1'b0;
  assign F2A_T_18_7 = 1'b0;
  assign F2A_T_1_0 = 1'b0;
  assign F2A_T_1_1 = 1'b0;
  assign F2A_T_1_10 = 1'b0;
  assign F2A_T_1_11 = 1'b0;
  assign F2A_T_1_2 = 1'b0;
  assign F2A_T_1_3 = 1'b0;
  assign F2A_T_1_4 = 1'b0;
  assign F2A_T_1_5 = 1'b0;
  assign F2A_T_1_6 = 1'b0;
  assign F2A_T_1_7 = 1'b0;
  assign F2A_T_1_8 = 1'b0;
  assign F2A_T_1_9 = 1'b0;
  assign F2A_T_23_11 = 1'b0;
  assign F2A_T_24_0 = 1'b0;
  assign F2A_T_24_1 = 1'b0;
  assign F2A_T_24_10 = 1'b0;
  assign F2A_T_24_11 = 1'b0;
  assign F2A_T_24_12 = 1'b0;
  assign F2A_T_24_13 = 1'b0;
  assign F2A_T_24_14 = 1'b0;
  assign F2A_T_24_15 = 1'b0;
  assign F2A_T_24_2 = 1'b0;
  assign F2A_T_24_3 = 1'b0;
  assign F2A_T_24_4 = 1'b0;
  assign F2A_T_24_5 = 1'b0;
  assign F2A_T_24_6 = 1'b0;
  assign F2A_T_24_7 = 1'b0;
  assign F2A_T_24_8 = 1'b0;
  assign F2A_T_24_9 = 1'b0;
  assign F2A_T_28_10 = 1'b0;
  assign F2A_T_28_11 = 1'b0;
  assign F2A_T_28_12 = 1'b0;
  assign F2A_T_28_13 = 1'b0;
  assign F2A_T_28_14 = 1'b0;
  assign F2A_T_28_5 = 1'b0;
  assign F2A_T_28_6 = 1'b0;
  assign F2A_T_28_7 = 1'b0;
  assign F2A_T_28_8 = 1'b0;
  assign F2A_T_28_9 = 1'b0;
  assign F2A_T_30_0 = 1'b0;
  assign F2A_T_30_1 = 1'b0;
  assign F2A_T_30_10 = 1'b0;
  assign F2A_T_30_11 = 1'b0;
  assign F2A_T_30_12 = 1'b0;
  assign F2A_T_30_13 = 1'b0;
  assign F2A_T_30_14 = 1'b0;
  assign F2A_T_30_15 = 1'b0;
  assign F2A_T_30_16 = 1'b0;
  assign F2A_T_30_17 = 1'b0;
  assign F2A_T_30_2 = 1'b0;
  assign F2A_T_30_3 = 1'b0;
  assign F2A_T_30_4 = 1'b0;
  assign F2A_T_30_5 = 1'b0;
  assign F2A_T_30_6 = 1'b0;
  assign F2A_T_30_7 = 1'b0;
  assign F2A_T_30_8 = 1'b0;
  assign F2A_T_30_9 = 1'b0;
  assign F2A_T_31_0 = 1'b0;
  assign F2A_T_31_1 = 1'b0;
  assign F2A_T_31_10 = 1'b0;
  assign F2A_T_31_11 = 1'b0;
  assign F2A_T_31_2 = 1'b0;
  assign F2A_T_31_3 = 1'b0;
  assign F2A_T_31_4 = 1'b0;
  assign F2A_T_31_5 = 1'b0;
  assign F2A_T_31_6 = 1'b0;
  assign F2A_T_31_7 = 1'b0;
  assign F2A_T_31_8 = 1'b0;
  assign F2A_T_31_9 = 1'b0;
  assign F2A_T_32_0 = 1'b0;
  assign F2A_T_32_1 = 1'b0;
  assign F2A_T_32_10 = 1'b0;
  assign F2A_T_32_11 = 1'b0;
  assign F2A_T_32_12 = 1'b0;
  assign F2A_T_32_13 = 1'b0;
  assign F2A_T_32_14 = 1'b0;
  assign F2A_T_32_15 = 1'b0;
  assign F2A_T_32_16 = 1'b0;
  assign F2A_T_32_17 = 1'b0;
  assign F2A_T_32_2 = 1'b0;
  assign F2A_T_32_3 = 1'b0;
  assign F2A_T_32_4 = 1'b0;
  assign F2A_T_32_5 = 1'b0;
  assign F2A_T_32_6 = 1'b0;
  assign F2A_T_32_7 = 1'b0;
  assign F2A_T_32_8 = 1'b0;
  assign F2A_T_32_9 = 1'b0;
  assign F2Adef_B_10_0 = 1'b0;
  assign F2Adef_B_10_1 = 1'b0;
  assign F2Adef_B_10_2 = 1'b0;
  assign F2Adef_B_10_3 = 1'b0;
  assign F2Adef_B_10_4 = 1'b0;
  assign F2Adef_B_10_5 = 1'b0;
  assign F2Adef_B_10_6 = 1'b0;
  assign F2Adef_B_11_0 = 1'b0;
  assign F2Adef_B_11_1 = 1'b0;
  assign F2Adef_B_11_2 = 1'b0;
  assign F2Adef_B_11_3 = 1'b0;
  assign F2Adef_B_12_0 = 1'b0;
  assign F2Adef_B_12_1 = 1'b0;
  assign F2Adef_B_12_2 = 1'b0;
  assign F2Adef_B_12_3 = 1'b0;
  assign F2Adef_B_12_4 = 1'b0;
  assign F2Adef_B_12_5 = 1'b0;
  assign F2Adef_B_12_6 = 1'b0;
  assign F2Adef_B_13_1 = 1'b0;
  assign F2Adef_B_13_2 = 1'b0;
  assign F2Adef_B_13_3 = 1'b0;
  assign F2Adef_B_14_0 = 1'b0;
  assign F2Adef_B_14_1 = 1'b0;
  assign F2Adef_B_14_2 = 1'b0;
  assign F2Adef_B_14_3 = 1'b0;
  assign F2Adef_B_14_4 = 1'b0;
  assign F2Adef_B_14_5 = 1'b0;
  assign F2Adef_B_14_6 = 1'b0;
  assign F2Adef_B_15_0 = 1'b0;
  assign F2Adef_B_15_1 = 1'b0;
  assign F2Adef_B_15_2 = 1'b0;
  assign F2Adef_B_15_3 = 1'b0;
  assign F2Adef_B_16_0 = 1'b0;
  assign F2Adef_B_16_1 = 1'b0;
  assign F2Adef_B_16_2 = 1'b0;
  assign F2Adef_B_16_3 = 1'b0;
  assign F2Adef_B_16_4 = 1'b0;
  assign F2Adef_B_16_5 = 1'b0;
  assign F2Adef_B_16_6 = 1'b0;
  assign F2Adef_B_17_0 = 1'b0;
  assign F2Adef_B_17_1 = 1'b0;
  assign F2Adef_B_17_2 = 1'b0;
  assign F2Adef_B_17_3 = 1'b0;
  assign F2Adef_B_18_0 = 1'b0;
  assign F2Adef_B_18_1 = 1'b0;
  assign F2Adef_B_18_2 = 1'b0;
  assign F2Adef_B_18_3 = 1'b0;
  assign F2Adef_B_18_4 = 1'b0;
  assign F2Adef_B_18_5 = 1'b0;
  assign F2Adef_B_18_6 = 1'b0;
  assign F2Adef_B_19_0 = 1'b0;
  assign F2Adef_B_19_1 = 1'b0;
  assign F2Adef_B_19_2 = 1'b0;
  assign F2Adef_B_19_3 = 1'b0;
  assign F2Adef_B_1_0 = 1'b0;
  assign F2Adef_B_1_1 = 1'b0;
  assign F2Adef_B_1_2 = 1'b0;
  assign F2Adef_B_1_3 = 1'b0;
  assign F2Adef_B_20_0 = 1'b0;
  assign F2Adef_B_20_1 = 1'b0;
  assign F2Adef_B_20_2 = 1'b0;
  assign F2Adef_B_20_3 = 1'b0;
  assign F2Adef_B_20_4 = 1'b0;
  assign F2Adef_B_20_5 = 1'b0;
  assign F2Adef_B_20_6 = 1'b0;
  assign F2Adef_B_21_0 = 1'b0;
  assign F2Adef_B_21_1 = 1'b0;
  assign F2Adef_B_21_2 = 1'b0;
  assign F2Adef_B_21_3 = 1'b0;
  assign F2Adef_B_22_0 = 1'b0;
  assign F2Adef_B_22_1 = 1'b0;
  assign F2Adef_B_22_2 = 1'b0;
  assign F2Adef_B_22_3 = 1'b0;
  assign F2Adef_B_22_4 = 1'b0;
  assign F2Adef_B_22_5 = 1'b0;
  assign F2Adef_B_22_6 = 1'b0;
  assign F2Adef_B_23_0 = 1'b0;
  assign F2Adef_B_23_1 = 1'b0;
  assign F2Adef_B_23_2 = 1'b0;
  assign F2Adef_B_23_3 = 1'b0;
  assign F2Adef_B_24_0 = 1'b0;
  assign F2Adef_B_24_2 = 1'b0;
  assign F2Adef_B_24_3 = 1'b0;
  assign F2Adef_B_24_4 = 1'b0;
  assign F2Adef_B_24_5 = 1'b0;
  assign F2Adef_B_24_6 = 1'b0;
  assign F2Adef_B_25_0 = 1'b0;
  assign F2Adef_B_25_1 = 1'b0;
  assign F2Adef_B_25_2 = 1'b0;
  assign F2Adef_B_25_3 = 1'b0;
  assign F2Adef_B_26_0 = 1'b0;
  assign F2Adef_B_26_1 = 1'b0;
  assign F2Adef_B_26_2 = 1'b0;
  assign F2Adef_B_26_3 = 1'b0;
  assign F2Adef_B_26_4 = 1'b0;
  assign F2Adef_B_26_5 = 1'b0;
  assign F2Adef_B_26_6 = 1'b0;
  assign F2Adef_B_27_0 = 1'b0;
  assign F2Adef_B_27_1 = 1'b0;
  assign F2Adef_B_27_2 = 1'b0;
  assign F2Adef_B_27_3 = 1'b0;
  assign F2Adef_B_28_0 = 1'b0;
  assign F2Adef_B_28_1 = 1'b0;
  assign F2Adef_B_28_2 = 1'b0;
  assign F2Adef_B_28_3 = 1'b0;
  assign F2Adef_B_28_4 = 1'b0;
  assign F2Adef_B_28_5 = 1'b0;
  assign F2Adef_B_28_6 = 1'b0;
  assign F2Adef_B_29_0 = 1'b0;
  assign F2Adef_B_29_1 = 1'b0;
  assign F2Adef_B_29_2 = 1'b0;
  assign F2Adef_B_29_3 = 1'b0;
  assign F2Adef_B_2_0 = 1'b0;
  assign F2Adef_B_2_1 = 1'b0;
  assign F2Adef_B_2_2 = 1'b0;
  assign F2Adef_B_2_3 = 1'b0;
  assign F2Adef_B_2_4 = 1'b0;
  assign F2Adef_B_2_5 = 1'b0;
  assign F2Adef_B_2_6 = 1'b0;
  assign F2Adef_B_30_0 = 1'b0;
  assign F2Adef_B_30_1 = 1'b0;
  assign F2Adef_B_30_2 = 1'b0;
  assign F2Adef_B_30_3 = 1'b0;
  assign F2Adef_B_30_4 = 1'b0;
  assign F2Adef_B_30_5 = 1'b0;
  assign F2Adef_B_30_6 = 1'b0;
  assign F2Adef_B_31_0 = 1'b0;
  assign F2Adef_B_31_1 = 1'b0;
  assign F2Adef_B_31_2 = 1'b0;
  assign F2Adef_B_31_3 = 1'b0;
  assign F2Adef_B_32_0 = 1'b0;
  assign F2Adef_B_32_1 = 1'b0;
  assign F2Adef_B_32_2 = 1'b0;
  assign F2Adef_B_32_3 = 1'b0;
  assign F2Adef_B_32_4 = 1'b0;
  assign F2Adef_B_32_5 = 1'b0;
  assign F2Adef_B_32_6 = 1'b0;
  assign F2Adef_B_3_0 = 1'b0;
  assign F2Adef_B_3_1 = 1'b0;
  assign F2Adef_B_3_2 = 1'b0;
  assign F2Adef_B_3_3 = 1'b0;
  assign F2Adef_B_4_0 = 1'b0;
  assign F2Adef_B_4_1 = 1'b0;
  assign F2Adef_B_4_2 = 1'b0;
  assign F2Adef_B_4_3 = 1'b0;
  assign F2Adef_B_4_4 = 1'b0;
  assign F2Adef_B_4_5 = 1'b0;
  assign F2Adef_B_4_6 = 1'b0;
  assign F2Adef_B_5_0 = 1'b0;
  assign F2Adef_B_5_1 = 1'b0;
  assign F2Adef_B_5_2 = 1'b0;
  assign F2Adef_B_5_3 = 1'b0;
  assign F2Adef_B_6_0 = 1'b0;
  assign F2Adef_B_6_2 = 1'b0;
  assign F2Adef_B_6_3 = 1'b0;
  assign F2Adef_B_6_4 = 1'b0;
  assign F2Adef_B_6_5 = 1'b0;
  assign F2Adef_B_6_6 = 1'b0;
  assign F2Adef_B_7_0 = 1'b0;
  assign F2Adef_B_7_1 = 1'b0;
  assign F2Adef_B_7_2 = 1'b0;
  assign F2Adef_B_7_3 = 1'b0;
  assign F2Adef_B_8_0 = 1'b0;
  assign F2Adef_B_8_1 = 1'b0;
  assign F2Adef_B_8_2 = 1'b0;
  assign F2Adef_B_8_3 = 1'b0;
  assign F2Adef_B_8_4 = 1'b0;
  assign F2Adef_B_8_5 = 1'b0;
  assign F2Adef_B_8_6 = 1'b0;
  assign F2Adef_B_9_0 = 1'b0;
  assign F2Adef_B_9_1 = 1'b0;
  assign F2Adef_B_9_2 = 1'b0;
  assign F2Adef_B_9_3 = 1'b0;
  assign F2Adef_L_10_0 = 1'b0;
  assign F2Adef_L_10_1 = 1'b0;
  assign F2Adef_L_10_2 = 1'b0;
  assign F2Adef_L_10_3 = 1'b0;
  assign F2Adef_L_10_4 = 1'b0;
  assign F2Adef_L_10_5 = 1'b0;
  assign F2Adef_L_10_6 = 1'b0;
  assign F2Adef_L_11_0 = 1'b0;
  assign F2Adef_L_11_1 = 1'b0;
  assign F2Adef_L_11_2 = 1'b0;
  assign F2Adef_L_11_3 = 1'b0;
  assign F2Adef_L_12_0 = 1'b0;
  assign F2Adef_L_12_1 = 1'b0;
  assign F2Adef_L_12_2 = 1'b0;
  assign F2Adef_L_12_3 = 1'b0;
  assign F2Adef_L_12_4 = 1'b0;
  assign F2Adef_L_12_5 = 1'b0;
  assign F2Adef_L_12_6 = 1'b0;
  assign F2Adef_L_13_0 = 1'b0;
  assign F2Adef_L_13_1 = 1'b0;
  assign F2Adef_L_13_2 = 1'b0;
  assign F2Adef_L_13_3 = 1'b0;
  assign F2Adef_L_14_0 = 1'b0;
  assign F2Adef_L_14_1 = 1'b0;
  assign F2Adef_L_14_2 = 1'b0;
  assign F2Adef_L_14_3 = 1'b0;
  assign F2Adef_L_14_4 = 1'b0;
  assign F2Adef_L_14_5 = 1'b0;
  assign F2Adef_L_14_6 = 1'b0;
  assign F2Adef_L_15_0 = 1'b0;
  assign F2Adef_L_15_1 = 1'b0;
  assign F2Adef_L_15_2 = 1'b0;
  assign F2Adef_L_15_3 = 1'b0;
  assign F2Adef_L_16_0 = 1'b0;
  assign F2Adef_L_16_1 = 1'b0;
  assign F2Adef_L_16_2 = 1'b0;
  assign F2Adef_L_16_3 = 1'b0;
  assign F2Adef_L_16_4 = 1'b0;
  assign F2Adef_L_16_5 = 1'b0;
  assign F2Adef_L_16_6 = 1'b0;
  assign F2Adef_L_17_0 = 1'b0;
  assign F2Adef_L_17_1 = 1'b0;
  assign F2Adef_L_17_2 = 1'b0;
  assign F2Adef_L_17_3 = 1'b0;
  assign F2Adef_L_18_0 = 1'b0;
  assign F2Adef_L_18_1 = 1'b0;
  assign F2Adef_L_18_2 = 1'b0;
  assign F2Adef_L_18_3 = 1'b0;
  assign F2Adef_L_18_4 = 1'b0;
  assign F2Adef_L_18_5 = 1'b0;
  assign F2Adef_L_18_6 = 1'b0;
  assign F2Adef_L_19_0 = 1'b0;
  assign F2Adef_L_19_1 = 1'b0;
  assign F2Adef_L_19_2 = 1'b0;
  assign F2Adef_L_19_3 = 1'b0;
  assign F2Adef_L_1_0 = 1'b0;
  assign F2Adef_L_1_1 = 1'b0;
  assign F2Adef_L_1_2 = 1'b0;
  assign F2Adef_L_1_3 = 1'b0;
  assign F2Adef_L_20_0 = 1'b0;
  assign F2Adef_L_20_1 = 1'b0;
  assign F2Adef_L_20_2 = 1'b0;
  assign F2Adef_L_20_3 = 1'b0;
  assign F2Adef_L_20_4 = 1'b0;
  assign F2Adef_L_20_5 = 1'b0;
  assign F2Adef_L_20_6 = 1'b0;
  assign F2Adef_L_21_0 = 1'b0;
  assign F2Adef_L_21_1 = 1'b0;
  assign F2Adef_L_21_2 = 1'b0;
  assign F2Adef_L_21_3 = 1'b0;
  assign F2Adef_L_22_0 = 1'b0;
  assign F2Adef_L_22_1 = 1'b0;
  assign F2Adef_L_22_2 = 1'b0;
  assign F2Adef_L_22_3 = 1'b0;
  assign F2Adef_L_22_4 = 1'b0;
  assign F2Adef_L_22_5 = 1'b0;
  assign F2Adef_L_22_6 = 1'b0;
  assign F2Adef_L_23_0 = 1'b0;
  assign F2Adef_L_23_1 = 1'b0;
  assign F2Adef_L_23_2 = 1'b0;
  assign F2Adef_L_23_3 = 1'b0;
  assign F2Adef_L_24_0 = 1'b0;
  assign F2Adef_L_24_1 = 1'b0;
  assign F2Adef_L_24_2 = 1'b0;
  assign F2Adef_L_24_3 = 1'b0;
  assign F2Adef_L_24_4 = 1'b0;
  assign F2Adef_L_24_5 = 1'b0;
  assign F2Adef_L_24_6 = 1'b0;
  assign F2Adef_L_25_0 = 1'b0;
  assign F2Adef_L_25_1 = 1'b0;
  assign F2Adef_L_25_2 = 1'b0;
  assign F2Adef_L_25_3 = 1'b0;
  assign F2Adef_L_26_0 = 1'b0;
  assign F2Adef_L_26_1 = 1'b0;
  assign F2Adef_L_26_2 = 1'b0;
  assign F2Adef_L_26_3 = 1'b0;
  assign F2Adef_L_26_4 = 1'b0;
  assign F2Adef_L_26_5 = 1'b0;
  assign F2Adef_L_26_6 = 1'b0;
  assign F2Adef_L_27_0 = 1'b0;
  assign F2Adef_L_27_1 = 1'b0;
  assign F2Adef_L_27_2 = 1'b0;
  assign F2Adef_L_27_3 = 1'b0;
  assign F2Adef_L_28_0 = 1'b0;
  assign F2Adef_L_28_1 = 1'b0;
  assign F2Adef_L_28_2 = 1'b0;
  assign F2Adef_L_28_3 = 1'b0;
  assign F2Adef_L_28_4 = 1'b0;
  assign F2Adef_L_28_5 = 1'b0;
  assign F2Adef_L_28_6 = 1'b0;
  assign F2Adef_L_29_0 = 1'b0;
  assign F2Adef_L_29_1 = 1'b0;
  assign F2Adef_L_29_2 = 1'b0;
  assign F2Adef_L_29_3 = 1'b0;
  assign F2Adef_L_30_0 = 1'b0;
  assign F2Adef_L_30_1 = 1'b0;
  assign F2Adef_L_30_2 = 1'b0;
  assign F2Adef_L_30_3 = 1'b0;
  assign F2Adef_L_30_4 = 1'b0;
  assign F2Adef_L_30_5 = 1'b0;
  assign F2Adef_L_30_6 = 1'b0;
  assign F2Adef_L_31_0 = 1'b0;
  assign F2Adef_L_31_1 = 1'b0;
  assign F2Adef_L_31_2 = 1'b0;
  assign F2Adef_L_31_3 = 1'b0;
  assign F2Adef_L_32_0 = 1'b0;
  assign F2Adef_L_32_1 = 1'b0;
  assign F2Adef_L_32_2 = 1'b0;
  assign F2Adef_L_32_3 = 1'b0;
  assign F2Adef_L_32_4 = 1'b0;
  assign F2Adef_L_32_5 = 1'b0;
  assign F2Adef_L_32_6 = 1'b0;
  assign F2Adef_L_3_0 = 1'b0;
  assign F2Adef_L_3_1 = 1'b0;
  assign F2Adef_L_3_2 = 1'b0;
  assign F2Adef_L_3_3 = 1'b0;
  assign F2Adef_L_4_1 = 1'b0;
  assign F2Adef_L_4_2 = 1'b0;
  assign F2Adef_L_4_3 = 1'b0;
  assign F2Adef_L_4_4 = 1'b0;
  assign F2Adef_L_4_5 = 1'b0;
  assign F2Adef_L_4_6 = 1'b0;
  assign F2Adef_L_5_0 = 1'b0;
  assign F2Adef_L_5_1 = 1'b0;
  assign F2Adef_L_5_2 = 1'b0;
  assign F2Adef_L_5_3 = 1'b0;
  assign F2Adef_L_6_0 = 1'b0;
  assign F2Adef_L_6_1 = 1'b0;
  assign F2Adef_L_6_2 = 1'b0;
  assign F2Adef_L_6_3 = 1'b0;
  assign F2Adef_L_6_4 = 1'b0;
  assign F2Adef_L_6_5 = 1'b0;
  assign F2Adef_L_6_6 = 1'b0;
  assign F2Adef_L_7_0 = 1'b0;
  assign F2Adef_L_7_1 = 1'b0;
  assign F2Adef_L_7_2 = 1'b0;
  assign F2Adef_L_7_3 = 1'b0;
  assign F2Adef_L_8_0 = 1'b0;
  assign F2Adef_L_8_1 = 1'b0;
  assign F2Adef_L_8_2 = 1'b0;
  assign F2Adef_L_8_3 = 1'b0;
  assign F2Adef_L_8_4 = 1'b0;
  assign F2Adef_L_8_5 = 1'b0;
  assign F2Adef_L_8_6 = 1'b0;
  assign F2Adef_L_9_0 = 1'b0;
  assign F2Adef_L_9_1 = 1'b0;
  assign F2Adef_L_9_2 = 1'b0;
  assign F2Adef_L_9_3 = 1'b0;
  assign F2Adef_R_10_0 = 1'b0;
  assign F2Adef_R_10_1 = 1'b0;
  assign F2Adef_R_10_2 = 1'b0;
  assign F2Adef_R_10_3 = 1'b0;
  assign F2Adef_R_10_4 = 1'b0;
  assign F2Adef_R_10_5 = 1'b0;
  assign F2Adef_R_10_6 = 1'b0;
  assign F2Adef_R_11_0 = 1'b0;
  assign F2Adef_R_11_1 = 1'b0;
  assign F2Adef_R_11_2 = 1'b0;
  assign F2Adef_R_11_3 = 1'b0;
  assign F2Adef_R_12_0 = 1'b0;
  assign F2Adef_R_12_1 = 1'b0;
  assign F2Adef_R_12_2 = 1'b0;
  assign F2Adef_R_12_3 = 1'b0;
  assign F2Adef_R_12_4 = 1'b0;
  assign F2Adef_R_12_5 = 1'b0;
  assign F2Adef_R_12_6 = 1'b0;
  assign F2Adef_R_13_0 = 1'b0;
  assign F2Adef_R_13_1 = 1'b0;
  assign F2Adef_R_13_2 = 1'b0;
  assign F2Adef_R_13_3 = 1'b0;
  assign F2Adef_R_14_0 = 1'b0;
  assign F2Adef_R_14_1 = 1'b0;
  assign F2Adef_R_14_2 = 1'b0;
  assign F2Adef_R_14_3 = 1'b0;
  assign F2Adef_R_14_4 = 1'b0;
  assign F2Adef_R_14_5 = 1'b0;
  assign F2Adef_R_14_6 = 1'b0;
  assign F2Adef_R_15_0 = 1'b0;
  assign F2Adef_R_15_1 = 1'b0;
  assign F2Adef_R_15_2 = 1'b0;
  assign F2Adef_R_15_3 = 1'b0;
  assign F2Adef_R_16_0 = 1'b0;
  assign F2Adef_R_16_1 = 1'b0;
  assign F2Adef_R_16_2 = 1'b0;
  assign F2Adef_R_16_3 = 1'b0;
  assign F2Adef_R_16_4 = 1'b0;
  assign F2Adef_R_16_5 = 1'b0;
  assign F2Adef_R_16_6 = 1'b0;
  assign F2Adef_R_17_0 = 1'b0;
  assign F2Adef_R_17_1 = 1'b0;
  assign F2Adef_R_17_2 = 1'b0;
  assign F2Adef_R_17_3 = 1'b0;
  assign F2Adef_R_18_0 = 1'b0;
  assign F2Adef_R_18_1 = 1'b0;
  assign F2Adef_R_18_2 = 1'b0;
  assign F2Adef_R_18_3 = 1'b0;
  assign F2Adef_R_18_4 = 1'b0;
  assign F2Adef_R_18_5 = 1'b0;
  assign F2Adef_R_18_6 = 1'b0;
  assign F2Adef_R_19_0 = 1'b0;
  assign F2Adef_R_19_1 = 1'b0;
  assign F2Adef_R_19_2 = 1'b0;
  assign F2Adef_R_19_3 = 1'b0;
  assign F2Adef_R_1_0 = 1'b0;
  assign F2Adef_R_1_1 = 1'b0;
  assign F2Adef_R_1_2 = 1'b0;
  assign F2Adef_R_1_3 = 1'b0;
  assign F2Adef_R_20_0 = 1'b0;
  assign F2Adef_R_20_1 = 1'b0;
  assign F2Adef_R_20_2 = 1'b0;
  assign F2Adef_R_20_3 = 1'b0;
  assign F2Adef_R_20_4 = 1'b0;
  assign F2Adef_R_20_5 = 1'b0;
  assign F2Adef_R_20_6 = 1'b0;
  assign F2Adef_R_21_0 = 1'b0;
  assign F2Adef_R_21_1 = 1'b0;
  assign F2Adef_R_21_2 = 1'b0;
  assign F2Adef_R_21_3 = 1'b0;
  assign F2Adef_R_22_0 = 1'b0;
  assign F2Adef_R_22_1 = 1'b0;
  assign F2Adef_R_22_2 = 1'b0;
  assign F2Adef_R_22_3 = 1'b0;
  assign F2Adef_R_22_4 = 1'b0;
  assign F2Adef_R_22_5 = 1'b0;
  assign F2Adef_R_22_6 = 1'b0;
  assign F2Adef_R_23_0 = 1'b0;
  assign F2Adef_R_23_1 = 1'b0;
  assign F2Adef_R_23_2 = 1'b0;
  assign F2Adef_R_23_3 = 1'b0;
  assign F2Adef_R_24_0 = 1'b0;
  assign F2Adef_R_24_1 = 1'b0;
  assign F2Adef_R_24_2 = 1'b0;
  assign F2Adef_R_24_3 = 1'b0;
  assign F2Adef_R_24_4 = 1'b0;
  assign F2Adef_R_24_5 = 1'b0;
  assign F2Adef_R_24_6 = 1'b0;
  assign F2Adef_R_25_0 = 1'b0;
  assign F2Adef_R_25_1 = 1'b0;
  assign F2Adef_R_25_2 = 1'b0;
  assign F2Adef_R_25_3 = 1'b0;
  assign F2Adef_R_26_0 = 1'b0;
  assign F2Adef_R_26_1 = 1'b0;
  assign F2Adef_R_26_2 = 1'b0;
  assign F2Adef_R_26_3 = 1'b0;
  assign F2Adef_R_26_4 = 1'b0;
  assign F2Adef_R_26_5 = 1'b0;
  assign F2Adef_R_26_6 = 1'b0;
  assign F2Adef_R_27_0 = 1'b0;
  assign F2Adef_R_27_1 = 1'b0;
  assign F2Adef_R_27_2 = 1'b0;
  assign F2Adef_R_27_3 = 1'b0;
  assign F2Adef_R_28_0 = 1'b0;
  assign F2Adef_R_28_1 = 1'b0;
  assign F2Adef_R_28_2 = 1'b0;
  assign F2Adef_R_28_3 = 1'b0;
  assign F2Adef_R_28_4 = 1'b0;
  assign F2Adef_R_28_5 = 1'b0;
  assign F2Adef_R_28_6 = 1'b0;
  assign F2Adef_R_29_0 = 1'b0;
  assign F2Adef_R_29_1 = 1'b0;
  assign F2Adef_R_29_2 = 1'b0;
  assign F2Adef_R_29_3 = 1'b0;
  assign F2Adef_R_2_0 = 1'b0;
  assign F2Adef_R_2_1 = 1'b0;
  assign F2Adef_R_2_2 = 1'b0;
  assign F2Adef_R_2_3 = 1'b0;
  assign F2Adef_R_2_4 = 1'b0;
  assign F2Adef_R_2_5 = 1'b0;
  assign F2Adef_R_2_6 = 1'b0;
  assign F2Adef_R_30_0 = 1'b0;
  assign F2Adef_R_30_1 = 1'b0;
  assign F2Adef_R_30_2 = 1'b0;
  assign F2Adef_R_30_3 = 1'b0;
  assign F2Adef_R_30_4 = 1'b0;
  assign F2Adef_R_30_5 = 1'b0;
  assign F2Adef_R_30_6 = 1'b0;
  assign F2Adef_R_31_0 = 1'b0;
  assign F2Adef_R_31_1 = 1'b0;
  assign F2Adef_R_31_2 = 1'b0;
  assign F2Adef_R_31_3 = 1'b0;
  assign F2Adef_R_32_0 = 1'b0;
  assign F2Adef_R_32_1 = 1'b0;
  assign F2Adef_R_32_2 = 1'b0;
  assign F2Adef_R_32_3 = 1'b0;
  assign F2Adef_R_32_4 = 1'b0;
  assign F2Adef_R_32_5 = 1'b0;
  assign F2Adef_R_32_6 = 1'b0;
  assign F2Adef_R_3_0 = 1'b0;
  assign F2Adef_R_3_1 = 1'b0;
  assign F2Adef_R_3_2 = 1'b0;
  assign F2Adef_R_3_3 = 1'b0;
  assign F2Adef_R_4_0 = 1'b0;
  assign F2Adef_R_4_1 = 1'b0;
  assign F2Adef_R_4_2 = 1'b0;
  assign F2Adef_R_4_3 = 1'b0;
  assign F2Adef_R_4_4 = 1'b0;
  assign F2Adef_R_4_5 = 1'b0;
  assign F2Adef_R_4_6 = 1'b0;
  assign F2Adef_R_5_0 = 1'b0;
  assign F2Adef_R_5_1 = 1'b0;
  assign F2Adef_R_5_2 = 1'b0;
  assign F2Adef_R_5_3 = 1'b0;
  assign F2Adef_R_6_0 = 1'b0;
  assign F2Adef_R_6_1 = 1'b0;
  assign F2Adef_R_6_2 = 1'b0;
  assign F2Adef_R_6_3 = 1'b0;
  assign F2Adef_R_6_4 = 1'b0;
  assign F2Adef_R_6_5 = 1'b0;
  assign F2Adef_R_6_6 = 1'b0;
  assign F2Adef_R_7_0 = 1'b0;
  assign F2Adef_R_7_1 = 1'b0;
  assign F2Adef_R_7_2 = 1'b0;
  assign F2Adef_R_7_3 = 1'b0;
  assign F2Adef_R_8_0 = 1'b0;
  assign F2Adef_R_8_1 = 1'b0;
  assign F2Adef_R_8_2 = 1'b0;
  assign F2Adef_R_8_3 = 1'b0;
  assign F2Adef_R_8_4 = 1'b0;
  assign F2Adef_R_8_5 = 1'b0;
  assign F2Adef_R_8_6 = 1'b0;
  assign F2Adef_R_9_0 = 1'b0;
  assign F2Adef_R_9_1 = 1'b0;
  assign F2Adef_R_9_2 = 1'b0;
  assign F2Adef_R_9_3 = 1'b0;
  assign F2Adef_T_10_0 = 1'b0;
  assign F2Adef_T_10_1 = 1'b0;
  assign F2Adef_T_10_2 = 1'b0;
  assign F2Adef_T_10_3 = 1'b0;
  assign F2Adef_T_10_4 = 1'b0;
  assign F2Adef_T_10_5 = 1'b0;
  assign F2Adef_T_10_6 = 1'b0;
  assign F2Adef_T_11_0 = 1'b0;
  assign F2Adef_T_11_1 = 1'b0;
  assign F2Adef_T_11_2 = 1'b0;
  assign F2Adef_T_11_3 = 1'b0;
  assign F2Adef_T_12_0 = 1'b0;
  assign F2Adef_T_12_1 = 1'b0;
  assign F2Adef_T_12_2 = 1'b0;
  assign F2Adef_T_12_3 = 1'b0;
  assign F2Adef_T_12_4 = 1'b0;
  assign F2Adef_T_12_5 = 1'b0;
  assign F2Adef_T_12_6 = 1'b0;
  assign F2Adef_T_13_1 = 1'b0;
  assign F2Adef_T_13_2 = 1'b0;
  assign F2Adef_T_13_3 = 1'b0;
  assign F2Adef_T_14_0 = 1'b0;
  assign F2Adef_T_14_1 = 1'b0;
  assign F2Adef_T_14_2 = 1'b0;
  assign F2Adef_T_14_3 = 1'b0;
  assign F2Adef_T_14_4 = 1'b0;
  assign F2Adef_T_14_5 = 1'b0;
  assign F2Adef_T_14_6 = 1'b0;
  assign F2Adef_T_15_0 = 1'b0;
  assign F2Adef_T_15_1 = 1'b0;
  assign F2Adef_T_15_2 = 1'b0;
  assign F2Adef_T_15_3 = 1'b0;
  assign F2Adef_T_16_0 = 1'b0;
  assign F2Adef_T_16_1 = 1'b0;
  assign F2Adef_T_16_2 = 1'b0;
  assign F2Adef_T_16_3 = 1'b0;
  assign F2Adef_T_16_4 = 1'b0;
  assign F2Adef_T_16_5 = 1'b0;
  assign F2Adef_T_16_6 = 1'b0;
  assign F2Adef_T_17_0 = 1'b0;
  assign F2Adef_T_17_1 = 1'b0;
  assign F2Adef_T_17_2 = 1'b0;
  assign F2Adef_T_17_3 = 1'b0;
  assign F2Adef_T_18_0 = 1'b0;
  assign F2Adef_T_18_1 = 1'b0;
  assign F2Adef_T_18_2 = 1'b0;
  assign F2Adef_T_18_3 = 1'b0;
  assign F2Adef_T_18_4 = 1'b0;
  assign F2Adef_T_18_5 = 1'b0;
  assign F2Adef_T_18_6 = 1'b0;
  assign F2Adef_T_19_0 = 1'b0;
  assign F2Adef_T_19_1 = 1'b0;
  assign F2Adef_T_19_2 = 1'b0;
  assign F2Adef_T_19_3 = 1'b0;
  assign F2Adef_T_1_0 = 1'b0;
  assign F2Adef_T_1_1 = 1'b0;
  assign F2Adef_T_1_2 = 1'b0;
  assign F2Adef_T_1_3 = 1'b0;
  assign F2Adef_T_20_0 = 1'b0;
  assign F2Adef_T_20_1 = 1'b0;
  assign F2Adef_T_20_2 = 1'b0;
  assign F2Adef_T_20_3 = 1'b0;
  assign F2Adef_T_20_4 = 1'b0;
  assign F2Adef_T_20_5 = 1'b0;
  assign F2Adef_T_20_6 = 1'b0;
  assign F2Adef_T_21_0 = 1'b0;
  assign F2Adef_T_21_1 = 1'b0;
  assign F2Adef_T_21_2 = 1'b0;
  assign F2Adef_T_21_3 = 1'b0;
  assign F2Adef_T_22_0 = 1'b0;
  assign F2Adef_T_22_1 = 1'b0;
  assign F2Adef_T_22_2 = 1'b0;
  assign F2Adef_T_22_3 = 1'b0;
  assign F2Adef_T_22_4 = 1'b0;
  assign F2Adef_T_22_5 = 1'b0;
  assign F2Adef_T_22_6 = 1'b0;
  assign F2Adef_T_23_0 = 1'b0;
  assign F2Adef_T_23_1 = 1'b0;
  assign F2Adef_T_23_2 = 1'b0;
  assign F2Adef_T_23_3 = 1'b0;
  assign F2Adef_T_24_1 = 1'b0;
  assign F2Adef_T_24_2 = 1'b0;
  assign F2Adef_T_24_3 = 1'b0;
  assign F2Adef_T_24_4 = 1'b0;
  assign F2Adef_T_24_5 = 1'b0;
  assign F2Adef_T_24_6 = 1'b0;
  assign F2Adef_T_25_0 = 1'b0;
  assign F2Adef_T_25_1 = 1'b0;
  assign F2Adef_T_25_2 = 1'b0;
  assign F2Adef_T_25_3 = 1'b0;
  assign F2Adef_T_26_0 = 1'b0;
  assign F2Adef_T_26_1 = 1'b0;
  assign F2Adef_T_26_2 = 1'b0;
  assign F2Adef_T_26_3 = 1'b0;
  assign F2Adef_T_26_4 = 1'b0;
  assign F2Adef_T_26_5 = 1'b0;
  assign F2Adef_T_26_6 = 1'b0;
  assign F2Adef_T_27_0 = 1'b0;
  assign F2Adef_T_27_1 = 1'b0;
  assign F2Adef_T_27_2 = 1'b0;
  assign F2Adef_T_27_3 = 1'b0;
  assign F2Adef_T_28_0 = 1'b0;
  assign F2Adef_T_28_1 = 1'b0;
  assign F2Adef_T_28_2 = 1'b0;
  assign F2Adef_T_28_3 = 1'b0;
  assign F2Adef_T_28_4 = 1'b0;
  assign F2Adef_T_28_5 = 1'b0;
  assign F2Adef_T_28_6 = 1'b0;
  assign F2Adef_T_29_0 = 1'b0;
  assign F2Adef_T_29_1 = 1'b0;
  assign F2Adef_T_29_2 = 1'b0;
  assign F2Adef_T_29_3 = 1'b0;
  assign F2Adef_T_2_0 = 1'b0;
  assign F2Adef_T_2_1 = 1'b0;
  assign F2Adef_T_2_2 = 1'b0;
  assign F2Adef_T_2_3 = 1'b0;
  assign F2Adef_T_2_4 = 1'b0;
  assign F2Adef_T_2_5 = 1'b0;
  assign F2Adef_T_2_6 = 1'b0;
  assign F2Adef_T_30_0 = 1'b0;
  assign F2Adef_T_30_1 = 1'b0;
  assign F2Adef_T_30_2 = 1'b0;
  assign F2Adef_T_30_3 = 1'b0;
  assign F2Adef_T_30_4 = 1'b0;
  assign F2Adef_T_30_5 = 1'b0;
  assign F2Adef_T_30_6 = 1'b0;
  assign F2Adef_T_31_0 = 1'b0;
  assign F2Adef_T_31_1 = 1'b0;
  assign F2Adef_T_31_2 = 1'b0;
  assign F2Adef_T_31_3 = 1'b0;
  assign F2Adef_T_32_0 = 1'b0;
  assign F2Adef_T_32_1 = 1'b0;
  assign F2Adef_T_32_2 = 1'b0;
  assign F2Adef_T_32_3 = 1'b0;
  assign F2Adef_T_32_4 = 1'b0;
  assign F2Adef_T_32_5 = 1'b0;
  assign F2Adef_T_32_6 = 1'b0;
  assign F2Adef_T_3_0 = 1'b0;
  assign F2Adef_T_3_1 = 1'b0;
  assign F2Adef_T_3_2 = 1'b0;
  assign F2Adef_T_3_3 = 1'b0;
  assign F2Adef_T_4_0 = 1'b0;
  assign F2Adef_T_4_1 = 1'b0;
  assign F2Adef_T_4_2 = 1'b0;
  assign F2Adef_T_4_3 = 1'b0;
  assign F2Adef_T_4_4 = 1'b0;
  assign F2Adef_T_4_5 = 1'b0;
  assign F2Adef_T_4_6 = 1'b0;
  assign F2Adef_T_5_0 = 1'b0;
  assign F2Adef_T_5_1 = 1'b0;
  assign F2Adef_T_5_2 = 1'b0;
  assign F2Adef_T_5_3 = 1'b0;
  assign F2Adef_T_6_0 = 1'b0;
  assign F2Adef_T_6_2 = 1'b0;
  assign F2Adef_T_6_3 = 1'b0;
  assign F2Adef_T_6_4 = 1'b0;
  assign F2Adef_T_6_5 = 1'b0;
  assign F2Adef_T_6_6 = 1'b0;
  assign F2Adef_T_7_0 = 1'b0;
  assign F2Adef_T_7_1 = 1'b0;
  assign F2Adef_T_7_2 = 1'b0;
  assign F2Adef_T_7_3 = 1'b0;
  assign F2Adef_T_8_0 = 1'b0;
  assign F2Adef_T_8_1 = 1'b0;
  assign F2Adef_T_8_2 = 1'b0;
  assign F2Adef_T_8_3 = 1'b0;
  assign F2Adef_T_8_4 = 1'b0;
  assign F2Adef_T_8_5 = 1'b0;
  assign F2Adef_T_8_6 = 1'b0;
  assign F2Adef_T_9_0 = 1'b0;
  assign F2Adef_T_9_1 = 1'b0;
  assign F2Adef_T_9_2 = 1'b0;
  assign F2Adef_T_9_3 = 1'b0;
  assign F2Areg_B_11_0 = 1'b0;
  assign F2Areg_B_11_1 = 1'b0;
  assign F2Areg_B_13_0 = 1'b0;
  assign F2Areg_B_13_1 = 1'b0;
  assign F2Areg_B_15_0 = 1'b0;
  assign F2Areg_B_15_1 = 1'b0;
  assign F2Areg_B_17_0 = 1'b0;
  assign F2Areg_B_17_1 = 1'b0;
  assign F2Areg_B_19_0 = 1'b0;
  assign F2Areg_B_19_1 = 1'b0;
  assign F2Areg_B_1_0 = 1'b0;
  assign F2Areg_B_1_1 = 1'b0;
  assign F2Areg_B_21_0 = 1'b0;
  assign F2Areg_B_21_1 = 1'b0;
  assign F2Areg_B_23_0 = 1'b0;
  assign F2Areg_B_23_1 = 1'b0;
  assign F2Areg_B_25_0 = 1'b0;
  assign F2Areg_B_25_1 = 1'b0;
  assign F2Areg_B_27_0 = 1'b0;
  assign F2Areg_B_27_1 = 1'b0;
  assign F2Areg_B_29_0 = 1'b0;
  assign F2Areg_B_29_1 = 1'b0;
  assign F2Areg_B_31_0 = 1'b0;
  assign F2Areg_B_31_1 = 1'b0;
  assign F2Areg_B_3_0 = 1'b0;
  assign F2Areg_B_3_1 = 1'b0;
  assign F2Areg_B_5_0 = 1'b0;
  assign F2Areg_B_5_1 = 1'b0;
  assign F2Areg_B_7_0 = 1'b0;
  assign F2Areg_B_7_1 = 1'b0;
  assign F2Areg_B_9_0 = 1'b0;
  assign F2Areg_B_9_1 = 1'b0;
  assign F2Areg_L_11_0 = 1'b0;
  assign F2Areg_L_11_1 = 1'b0;
  assign F2Areg_L_13_0 = 1'b0;
  assign F2Areg_L_13_1 = 1'b0;
  assign F2Areg_L_15_0 = 1'b0;
  assign F2Areg_L_15_1 = 1'b0;
  assign F2Areg_L_17_0 = 1'b0;
  assign F2Areg_L_17_1 = 1'b0;
  assign F2Areg_L_19_0 = 1'b0;
  assign F2Areg_L_19_1 = 1'b0;
  assign F2Areg_L_1_0 = 1'b0;
  assign F2Areg_L_1_1 = 1'b0;
  assign F2Areg_L_21_0 = 1'b0;
  assign F2Areg_L_21_1 = 1'b0;
  assign F2Areg_L_23_0 = 1'b0;
  assign F2Areg_L_23_1 = 1'b0;
  assign F2Areg_L_25_0 = 1'b0;
  assign F2Areg_L_25_1 = 1'b0;
  assign F2Areg_L_27_0 = 1'b0;
  assign F2Areg_L_27_1 = 1'b0;
  assign F2Areg_L_29_0 = 1'b0;
  assign F2Areg_L_29_1 = 1'b0;
  assign F2Areg_L_31_0 = 1'b0;
  assign F2Areg_L_31_1 = 1'b0;
  assign F2Areg_L_3_0 = 1'b0;
  assign F2Areg_L_3_1 = 1'b0;
  assign F2Areg_L_5_0 = 1'b0;
  assign F2Areg_L_5_1 = 1'b0;
  assign F2Areg_L_7_0 = 1'b0;
  assign F2Areg_L_7_1 = 1'b0;
  assign F2Areg_L_9_0 = 1'b0;
  assign F2Areg_L_9_1 = 1'b0;
  assign F2Areg_R_11_0 = 1'b0;
  assign F2Areg_R_11_1 = 1'b0;
  assign F2Areg_R_13_0 = 1'b0;
  assign F2Areg_R_13_1 = 1'b0;
  assign F2Areg_R_15_0 = 1'b0;
  assign F2Areg_R_15_1 = 1'b0;
  assign F2Areg_R_17_0 = 1'b0;
  assign F2Areg_R_17_1 = 1'b0;
  assign F2Areg_R_19_0 = 1'b0;
  assign F2Areg_R_19_1 = 1'b0;
  assign F2Areg_R_1_0 = 1'b0;
  assign F2Areg_R_1_1 = 1'b0;
  assign F2Areg_R_21_0 = 1'b0;
  assign F2Areg_R_21_1 = 1'b0;
  assign F2Areg_R_23_0 = 1'b0;
  assign F2Areg_R_23_1 = 1'b0;
  assign F2Areg_R_25_0 = 1'b0;
  assign F2Areg_R_25_1 = 1'b0;
  assign F2Areg_R_27_0 = 1'b0;
  assign F2Areg_R_27_1 = 1'b0;
  assign F2Areg_R_29_0 = 1'b0;
  assign F2Areg_R_29_1 = 1'b0;
  assign F2Areg_R_31_0 = 1'b0;
  assign F2Areg_R_31_1 = 1'b0;
  assign F2Areg_R_3_0 = 1'b0;
  assign F2Areg_R_3_1 = 1'b0;
  assign F2Areg_R_5_0 = 1'b0;
  assign F2Areg_R_5_1 = 1'b0;
  assign F2Areg_R_7_0 = 1'b0;
  assign F2Areg_R_7_1 = 1'b0;
  assign F2Areg_R_9_0 = 1'b0;
  assign F2Areg_R_9_1 = 1'b0;
  assign F2Areg_T_11_0 = 1'b0;
  assign F2Areg_T_11_1 = 1'b0;
  assign F2Areg_T_13_0 = 1'b0;
  assign F2Areg_T_13_1 = 1'b0;
  assign F2Areg_T_15_0 = 1'b0;
  assign F2Areg_T_15_1 = 1'b0;
  assign F2Areg_T_17_0 = 1'b0;
  assign F2Areg_T_17_1 = 1'b0;
  assign F2Areg_T_19_0 = 1'b0;
  assign F2Areg_T_19_1 = 1'b0;
  assign F2Areg_T_1_0 = 1'b0;
  assign F2Areg_T_1_1 = 1'b0;
  assign F2Areg_T_21_0 = 1'b0;
  assign F2Areg_T_21_1 = 1'b0;
  assign F2Areg_T_23_0 = 1'b0;
  assign F2Areg_T_23_1 = 1'b0;
  assign F2Areg_T_25_0 = 1'b0;
  assign F2Areg_T_25_1 = 1'b0;
  assign F2Areg_T_27_0 = 1'b0;
  assign F2Areg_T_27_1 = 1'b0;
  assign F2Areg_T_29_0 = 1'b0;
  assign F2Areg_T_29_1 = 1'b0;
  assign F2Areg_T_31_0 = 1'b0;
  assign F2Areg_T_31_1 = 1'b0;
  assign F2Areg_T_3_0 = 1'b0;
  assign F2Areg_T_3_1 = 1'b0;
  assign F2Areg_T_5_0 = 1'b0;
  assign F2Areg_T_5_1 = 1'b0;
  assign F2Areg_T_7_0 = 1'b0;
  assign F2Areg_T_7_1 = 1'b0;
  assign F2Areg_T_9_0 = 1'b0;
  assign F2Areg_T_9_1 = 1'b0;
endmodule
