
//--------------------------------------------------------------------------------//
//--										--//
//-- QuickLogic confidential 2016     					--// 
//--										--//
//-- File name 		: qf_rwhwsc.sv					--//	
//-- Create time 	: Fri Jul 15 14:53:54 2016				--// 
//-- Owner		: jcheng 					--//
//-- 										--//
//-- Function Description :							--//
//--										--//
//--										--//
//-- Modification 	 							--//
//-- 1. 									--//
//-- Date 		:							--//
//-- Owner 		:							--//
//-- Change(s) 		:							--//
//--										--//
//--										--//
//--										--//
//--------------------------------------------------------------------------------//

module qf_rwhwsc 
#(
parameter               PAR_BIT_WIDTH 		= 10 ,
parameter               PAR_DEFAULT_VALUE 	= 10'h000 
)
(
        //------------------------------------------------------------------------//
        //-- INPUT PORT                                                         --//
        //------------------------------------------------------------------------//
        	//----------------------------------------------------------------//
        	//-- CLK							--//
        	//----------------------------------------------------------------//
input logic				sys_clk ,
input logic				sys_rst_n ,
input logic [PAR_BIT_WIDTH -1 :0]       wrdata ,
input logic             		wr_en ,
input logic				hw_wr_en ,
input logic [PAR_BIT_WIDTH -1 :0]       hw_wrdata ,
        //------------------------------------------------------------------------//
        //-- OUTPUT PORT                                                        --//
        //------------------------------------------------------------------------//
output logic [PAR_BIT_WIDTH -1 :0]      rddata 
);
        //------------------------------------------------------------------------//
        //-- Declare Time Unit                                                  --//
        //------------------------------------------------------------------------//
timeunit                1ns;
timeprecision           100ps ;

        //------------------------------------------------------------------------//
        //-- Local Parameter                                                    --//
        //------------------------------------------------------------------------//
localparam              PAR_DLY = 1'b1 ;

        //------------------------------------------------------------------------//
        //-- Wire/Flops                                                         --//
        //------------------------------------------------------------------------//
logic [PAR_BIT_WIDTH - 1 :0]            data_cs ;
logic [PAR_BIT_WIDTH - 1 :0]            data_ns ;

//--------------------------------------------------------------------------------//
//-- Start Functional Description                                               --//
//--------------------------------------------------------------------------------//
        //------------------------------------------------------------------------//
        //--                                                                    --//
        //------------------------------------------------------------------------//
assign rddata = data_cs ;

        //------------------------------------------------------------------------//
        //-- SYNC                                                               --//
        //------------------------------------------------------------------------//
always_ff @ ( posedge sys_clk or negedge sys_rst_n )
begin
  if ( sys_rst_n == 1'b0 )
    begin
        data_cs <= #PAR_DLY PAR_DEFAULT_VALUE ;
    end
  else
    begin
        data_cs <= #PAR_DLY data_ns  ;
    end
end
        //------------------------------------------------------------------------//
        //-- COMB                                                               --//
        //------------------------------------------------------------------------//
always_comb
begin
  if ( hw_wr_en == 1'b1 )
    begin
      data_ns = hw_wrdata ;
    end
  else if ( wr_en == 1'b1 )
    begin
      data_ns = wrdata   ;
    end
  else 
    begin
      data_ns = data_cs  ;
    end
end
//--------------------------------------------------------------------------------//
//-- END                                                                        --//
//--------------------------------------------------------------------------------//
endmodule
