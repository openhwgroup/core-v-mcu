//Version : AU 1.3.0.PreRelease Oct 15 2020

module A2_design (
    input [5:0] CLK,
    input [3:0] RESET,

    input [31:0] m0_oper0_rdata,
    input [31:0] m0_m0_dataout,
    input [31:0] m0_coef_rdata,
    input [31:0] m0_m1_dataout,
    input [31:0] m0_oper1_rdata,
    input [31:0] m1_oper0_rdata,
    input [31:0] m1_m0_dataout,
    input [31:0] m1_coef_rdata,
    input [31:0] m1_m1_dataout,
    input [31:0] m1_oper1_rdata,

    input [79:0] fpgaio_in,
    input [31:0] lint_WDATA,
    input [19:0] lint_ADDR,
    input        lint_REQ,
    input        lint_WEN,
    input [ 3:0] lint_BE,
    input [31:0] control_in,

    input [31:0] tcdm_rdata_p0,
    input [31:0] tcdm_rdata_p1,
    input [31:0] tcdm_rdata_p2,
    input [31:0] tcdm_rdata_p3,

    input               tcdm_valid_p0,
    input               tcdm_gnt_p0,
    input               tcdm_fmo_p0,
    input               tcdm_valid_p1,
    input               tcdm_gnt_p1,
    input               tcdm_fmo_p1,
    input               tcdm_valid_p2,
    input               tcdm_gnt_p2,
    input               tcdm_fmo_p2,
    input               tcdm_valid_p3,
    input               tcdm_gnt_p3,
    input               tcdm_fmo_p3,
    input  logic [ 3:0] FB_SPE_IN,
    output logic [ 3:0] FB_SPE_OUT,
    inout  logic        NB,
    inout  logic        PB,
    input  logic        MLATCH,
    input  logic        POR,
    input  logic        STM,
    input  logic [ 5:0] M,
    input  logic [31:0] fcb_bl_din,
    output logic [31:0] fcb_bl_dout,
    input  logic [15:0] fcb_bl_pwrgate,
    input  logic        fcb_blclk,
    input  logic        fcb_cload_din_sel,
    input  logic        fcb_din_int_l_only,
    input  logic        fcb_din_int_r_only,
    input  logic        fcb_din_slc_tb_int,
    input  logic        fcb_fb_iso_enb,
    input  logic [15:0] fcb_iso_en,
    input  logic        fcb_pchg_b,
    input  logic [15:0] fcb_pi_pwr,
    output logic        fcb_pif_en,
    input  logic [15:0] fcb_prog,
    input  logic        fcb_prog_ifx,
    input  logic        fcb_pwr_gate,
    input  logic        fcb_re,
    input  logic [15:0] fcb_vlp_clkdis,
    input  logic        fcb_vlp_clkdis_ifx,
    input  logic [15:0] fcb_vlp_pwrdis,
    input  logic        fcb_vlp_pwrdis_ifx,
    input  logic [15:0] fcb_vlp_srdis,
    input  logic        fcb_vlp_srdis_ifx,
    input  logic        fcb_we,
    input  logic        fcb_we_int,
    input  logic [ 2:0] fcb_wl_cload_sel,
    input  logic [ 5:0] fcb_wl_din,
    input  logic        fcb_wl_en,
    input  logic        fcb_wl_int_din_sel,
    input  logic [ 7:0] fcb_wl_pwrgate,
    input  logic        fcb_wl_resetb,
    input  logic [15:0] fcb_wl_sel,
    input  logic        fcb_wl_sel_tb_int,
    input  logic        fcb_wlclk,

    input  logic        fcb_fb_cfg_done,
    output       [31:0] m0_m0_oper_in,
    output              m0_m0_osel,
    output       [31:0] m0_m0_coef_in,
    output              m0_m0_csel,
    output       [ 1:0] m0_m0_mode,
    output       [ 5:0] m0_m0_outsel,
    output              m0_m0_clk,
    output              m0_m0_reset,
    output              m0_m0_clken,
    output              m0_m0_clr,
    output              m0_m0_sat,
    output              m0_m0_rnd,
    output              m0_m0_tc,

    output [31:0] m0_m1_oper_in,
    output        m0_m1_osel,
    output [31:0] m0_m1_coef_in,
    output        m0_m1_csel,
    output [ 1:0] m0_m1_mode,
    output [ 5:0] m0_m1_outsel,
    output        m0_m1_clk,
    output        m0_m1_reset,
    output        m0_m1_clken,
    output        m0_m1_clr,
    output        m0_m1_sat,
    output        m0_m1_rnd,
    output        m0_m1_tc,

    output [31:0] m1_m0_oper_in,
    output        m1_m0_osel,
    output [31:0] m1_m0_coef_in,
    output        m1_m0_csel,
    output [ 1:0] m1_m0_mode,
    output [ 5:0] m1_m0_outsel,
    output        m1_m0_clk,
    output        m1_m0_reset,
    output        m1_m0_clken,
    output        m1_m0_clr,
    output        m1_m0_sat,
    output        m1_m0_rnd,
    output        m1_m0_tc,

    output [31:0] m1_m1_oper_in,
    output        m1_m1_osel,
    output [31:0] m1_m1_coef_in,
    output        m1_m1_csel,
    output [ 1:0] m1_m1_mode,
    output [ 5:0] m1_m1_outsel,
    output        m1_m1_clk,
    output        m1_m1_reset,
    output        m1_m1_clken,
    output        m1_m1_clr,
    output        m1_m1_sat,
    output        m1_m1_rnd,
    output        m1_m1_tc,

    output [31:0] m0_oper0_wdata,
    output [ 1:0] m0_oper0_rmode,
    output        m0_oper0_rclk,
    output [11:0] m0_oper0_raddr,
    output [11:0] m0_oper0_waddr,
    output [ 1:0] m0_oper0_wmode,
    output        m0_oper0_wclk,
    output        m0_oper0_we,
    output        m0_oper0_wdsel,
    output        m0_oper0_powerdn,

    output [31:0] m0_coef_wdata,
    output [ 1:0] m0_coef_rmode,
    output        m0_coef_rclk,
    output [11:0] m0_coef_raddr,
    output [11:0] m0_coef_waddr,

    output [1:0] m0_coef_wmode,
    output       m0_coef_wclk,
    output       m0_coef_we,
    output       m0_coef_wdsel,
    output       m0_coef_powerdn,

    output [31:0] m0_oper1_wdata,
    output [ 1:0] m0_oper1_rmode,
    output        m0_oper1_rclk,
    output [11:0] m0_oper1_raddr,
    output [11:0] m0_oper1_waddr,
    output [ 1:0] m0_oper1_wmode,
    output        m0_oper1_wclk,
    output        m0_oper1_we,
    output        m0_oper1_wdsel,
    output        m0_oper1_powerdn,

    output [31:0] m1_oper0_wdata,
    output [ 1:0] m1_oper0_rmode,
    output        m1_oper0_rclk,
    output [11:0] m1_oper0_raddr,
    output [11:0] m1_oper0_waddr,
    output [ 1:0] m1_oper0_wmode,
    output        m1_oper0_wclk,
    output        m1_oper0_we,
    output        m1_oper0_wdsel,
    output        m1_oper0_powerdn,

    output [31:0] m1_coef_wdata,
    output [ 1:0] m1_coef_rmode,
    output        m1_coef_rclk,
    output [11:0] m1_coef_raddr,
    output [11:0] m1_coef_waddr,
    output [ 1:0] m1_coef_wmode,
    output        m1_coef_wclk,
    output        m1_coef_we,
    output        m1_coef_wdsel,
    output        m1_coef_powerdn,

    output [31:0] m1_oper1_wdata,
    output [ 1:0] m1_oper1_rmode,
    output        m1_oper1_rclk,
    output [11:0] m1_oper1_raddr,
    output [11:0] m1_oper1_waddr,
    output [ 1:0] m1_oper1_wmode,
    output        m1_oper1_wclk,
    output        m1_oper1_we,
    output        m1_oper1_wdsel,
    output        m1_oper1_powerdn,

    output [79:0] fpgaio_out,
    output [79:0] fpgaio_oe,
    output [31:0] lint_RDATA,
    output        lint_clk,
    output        lint_VALID,
    output        lint_GNT,

    output [31:0] tcdm_wdata_p0,
    output [31:0] tcdm_wdata_p1,
    output [31:0] tcdm_wdata_p2,
    output [31:0] tcdm_wdata_p3,

    output [19:0] tcdm_addr_p0,
    output [19:0] tcdm_addr_p1,
    output [19:0] tcdm_addr_p2,
    output [19:0] tcdm_addr_p3,

    output       tcdm_wen_p0,
    tcdm_wen_p1,
    tcdm_wen_p2,
    tcdm_wen_p3,
    output       tcdm_clk_p0,
    output       tcdm_req_p0,
    output [3:0] tcdm_be_p0,

    output       tcdm_clk_p1,
    output       tcdm_req_p1,
    output [3:0] tcdm_be_p1,

    output       tcdm_clk_p2,
    output       tcdm_req_p2,
    output [3:0] tcdm_be_p2,

    output        tcdm_clk_p3,
    output        tcdm_req_p3,
    output [ 3:0] tcdm_be_p3,
    output [15:0] events_o,
    output [31:0] status_out,
    output [ 7:0] version,
    inout         VSSC,
    VDDC_FPGA
);


  // Gated clocks for SDC timing calculations

  wire m0_m0_clk_int, m0_m0_clk_def;
`ifndef FPGA
  pulp_clock_mux2 u1 (
      .clk0_i(m0_m0_clk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m0_m0_clk_def),
      .clk_o(m0_m0_clk)
  );
`else
  assign m0_m0_clk = m0_m0_clk_def ? CLK[0] : m0_m0_clk_int;
`endif
  wire m0_m1_clk_int, m0_m1_clk_def;
`ifndef FPGA
  pulp_clock_mux2 u2 (
      .clk0_i(m0_m1_clk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m0_m1_clk_def),
      .clk_o(m0_m1_clk)
  );
`else
  assign m0_m1_clk = m0_m1_clk_def ? CLK[0] : m0_m1_clk_int;
`endif

  wire m1_m0_clk_int, m1_m0_clk_def;
`ifndef FPGA
  pulp_clock_mux2 u3 (
      .clk0_i(m1_m0_clk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m1_m0_clk_def),
      .clk_o(m1_m0_clk)
  );
`else
  assign m1_m0_clk = m1_m0_clk_def ? CLK[0] : m1_m0_clk_int;
`endif

  wire m1_m1_clk_int, m1_m1_clk_def;
`ifndef FPGA
  pulp_clock_mux2 u4 (
      .clk0_i(m1_m1_clk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m1_m1_clk_def),
      .clk_o(m1_m1_clk)
  );
`else
  assign m1_m1_clk = m1_m1_clk_def ? CLK[0] : m1_m1_clk_int;
`endif

  wire m0_oper0_wclk_int, m0_oper0_wclk_def;
`ifndef FPGA
  pulp_clock_mux2 u5 (
      .clk0_i(m0_oper0_wclk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m0_oper0_wclk_def),
      .clk_o(m0_oper0_wclk)
  );
`else
  assign m0_oper0_wclk = m0_oper0_wclk_def ? CLK[0] : m0_oper0_wclk_int;
`endif

  wire m0_oper0_rclk_int, m0_oper0_rclk_def;
`ifndef FPGA
  pulp_clock_mux2 u6 (
      .clk0_i(m0_oper0_rclk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m0_oper0_rclk_def),
      .clk_o(m0_oper0_rclk)
  );
`else
  assign m0_oper0_rclk = m0_oper0_rclk_def ? CLK[0] : m0_oper0_rclk_int;
`endif

  wire m0_coef_wclk_int, m0_coef_wclk_def;
`ifndef FPGA
  pulp_clock_mux2 u7 (
      .clk0_i(m0_coef_wclk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m0_coef_wclk_def),
      .clk_o(m0_coef_wclk)
  );
`else
  assign m0_coef_wclk = m0_coef_wclk_def ? CLK[0] : m0_coef_wclk_int;
`endif

  wire m0_coef_rclk_int, m0_coef_rclk_def;
`ifndef FPGA
  pulp_clock_mux2 u8 (
      .clk0_i(m0_coef_rclk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m0_coef_rclk_def),
      .clk_o(m0_coef_rclk)
  );
`else
  assign m0_coef_rclk = m0_coef_rclk_def ? CLK[0] : m0_coef_rclk_int;
`endif

  wire m0_oper1_wclk_int, m0_oper1_wclk_def;
`ifndef FPGA
  pulp_clock_mux2 u9 (
      .clk0_i(m0_oper1_wclk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m0_oper1_wclk_def),
      .clk_o(m0_oper1_wclk)
  );
`else
  assign m0_oper1_wclk = m0_oper1_wclk_def ? CLK[0] : m0_oper1_wclk_int;
`endif

  wire m0_oper1_rclk_int, m0_oper1_rclk_def;
`ifndef FPGA
  pulp_clock_mux2 u10 (
      .clk0_i(m0_oper1_rclk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m0_oper1_rclk_def),
      .clk_o(m0_oper1_rclk)
  );
`else
  assign m0_oper1_rclk = m0_oper1_rclk_def ? CLK[0] : m0_oper1_rclk_int;
`endif

  wire m1_oper0_wclk_int, m1_oper0_wclk_def;
`ifndef FPGA
  pulp_clock_mux2 u11 (
      .clk0_i(m1_oper0_wclk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m1_oper0_wclk_def),
      .clk_o(m1_oper0_wclk)
  );
`else
  assign m1_oper0_wclk = m1_oper0_wclk_def ? CLK[0] : m1_oper0_wclk_int;
`endif

  wire m1_oper0_rclk_int, m1_oper0_rclk_def;
`ifndef FPGA
  pulp_clock_mux2 u12 (
      .clk0_i(m1_oper0_rclk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m1_oper0_rclk_def),
      .clk_o(m1_oper0_rclk)
  );
`else
  assign m1_oper0_rclk = m1_oper0_rclk_def ? CLK[0] : m1_oper0_rclk_int;
`endif

  wire m1_coef_wclk_int, m1_coef_wclk_def;
`ifndef FPGA
  pulp_clock_mux2 u13 (
      .clk0_i(m1_coef_wclk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m1_coef_wclk_def),
      .clk_o(m1_coef_wclk)
  );
`else
  assign m1_coef_wclk = m1_coef_wclk_def ? CLK[0] : m1_coef_wclk_int;
`endif

  wire m1_coef_rclk_int, m1_coef_rclk_def;
`ifndef FPGA
  pulp_clock_mux2 u14 (
      .clk0_i(m1_coef_rclk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m1_coef_rclk_def),
      .clk_o(m1_coef_rclk)
  );
`else
  assign m1_coef_rclk = m1_coef_rclk_def ? CLK[0] : m1_coef_rclk_int;
`endif

  wire m1_oper1_wclk_int, m1_oper1_wclk_def;
`ifndef FPGA
  pulp_clock_mux2 u15 (
      .clk0_i(m1_oper1_wclk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m1_oper1_wclk_def),
      .clk_o(m1_oper1_wclk)
  );
`else
  assign m1_oper1_wclk = m1_oper1_wclk_def ? CLK[0] : m1_oper1_wclk_int;
`endif

  wire m1_oper1_rclk_int, m1_oper1_rclk_def;

`ifndef FPGA
  pulp_clock_mux2 u16 (
      .clk0_i(m1_oper1_rclk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(m1_oper1_rclk_def),
      .clk_o(m1_oper1_rclk)
  );
`else
  assign m1_oper1_rclk = m1_oper1_rclk_def ? CLK[0] : m1_oper1_rclk_int;
`endif

  wire lint_clk_int, lint_clk_def;
`ifndef FPGA
  pulp_clock_mux2 u17 (
      .clk0_i(lint_clk_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(lint_clk_def),
      .clk_o(lint_clk)
  );
`else
  assign lint_clk = lint_clk_def ? CLK[0] : lint_clk_int;
`endif

  wire tcdm_clk_p0_int, tcdm_clk_p0_def;
`ifndef FPGA
  pulp_clock_mux2 u18 (
      .clk0_i(tcdm_clk_p0_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(tcdm_clk_p0_def),
      .clk_o(tcdm_clk_p0)
  );
`else
  assign tcdm_clk_p0 = tcdm_clk_p0_def ? CLK[0] : tcdm_clk_p0_int;
`endif

  wire tcdm_clk_p1_int, tcdm_clk_p1_def;
`ifndef FPGA
  pulp_clock_mux2 u19 (
      .clk0_i(tcdm_clk_p1_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(tcdm_clk_p1_def),
      .clk_o(tcdm_clk_p1)
  );
`else
  assign tcdm_clk_p1 = tcdm_clk_p1_def ? CLK[0] : tcdm_clk_p1_int;
`endif

  wire tcdm_clk_p2_int, tcdm_clk_p2_def;
`ifndef FPGA
  pulp_clock_mux2 u20 (
      .clk0_i(tcdm_clk_p2_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(tcdm_clk_p2_def),
      .clk_o(tcdm_clk_p2)
  );
`else
  assign tcdm_clk_p2 = tcdm_clk_p2_def ? CLK[0] : tcdm_clk_p2_int;
`endif

  wire tcdm_clk_p3_int, tcdm_clk_p3_def;
`ifndef FPGA
  pulp_clock_mux2 u21 (
      .clk0_i(tcdm_clk_p3_int),
      .clk1_i(CLK[0]),
      .clk_sel_i(tcdm_clk_p3_def),
      .clk_o(tcdm_clk_p3)
  );
`else
  assign tcdm_clk_p3 = tcdm_clk_p3_def ? CLK[0] : tcdm_clk_p3_int;
`endif




  //  ql737b_top A2 (
  QL_eFPGA_ArcticPro2_32X32_GF_22_Arnold2 A2 (
      //       .vddz(VDDC_FPGA),
      .A2F_CLK0(CLK[0]),
      .A2F_CLK1(CLK[1]),
      .A2F_CLK2(CLK[2]),
      .A2F_CLK3(CLK[3]),
      .A2F_CLK4(CLK[4]),
      .A2F_CLK5(CLK[5]),
      .A2F_B_10_0(m1_m0_dataout[11]),
      .A2F_B_10_1(m1_m0_dataout[10]),
      .A2F_B_10_2(m1_m0_dataout[9]),
      .A2F_B_10_3(m1_m0_dataout[8]),
      .A2F_B_10_4(m1_m0_dataout[7]),
      .A2F_B_10_5(m1_m0_dataout[6]),
      .A2F_B_10_6(m1_m0_dataout[5]),
      .A2F_B_10_7(m1_m0_dataout[4]),
      .A2F_B_11_0(m1_m0_dataout[3]),
      .A2F_B_11_1(m1_m0_dataout[2]),
      .A2F_B_11_2(m1_m0_dataout[1]),
      .A2F_B_11_3(m1_m0_dataout[0]),
      .A2F_B_11_4(m1_coef_rdata[31]),
      .A2F_B_11_5(m1_coef_rdata[30]),
      .A2F_B_12_0(m1_coef_rdata[29]),
      .A2F_B_12_1(m1_coef_rdata[28]),
      .A2F_B_12_2(m1_coef_rdata[27]),
      .A2F_B_12_3(m1_coef_rdata[26]),
      .A2F_B_12_4(m1_coef_rdata[25]),
      .A2F_B_12_5(m1_coef_rdata[24]),
      .A2F_B_12_6(m1_coef_rdata[23]),
      .A2F_B_12_7(m1_coef_rdata[22]),
      .A2F_B_13_0(m1_coef_rdata[21]),
      .A2F_B_13_1(m1_coef_rdata[20]),
      .A2F_B_13_2(m1_coef_rdata[19]),
      .A2F_B_13_3(m1_coef_rdata[18]),
      .A2F_B_13_4(m1_coef_rdata[17]),
      .A2F_B_13_5(m1_coef_rdata[16]),
      .A2F_B_14_0(m1_coef_rdata[15]),
      .A2F_B_14_1(m1_coef_rdata[14]),
      .A2F_B_14_2(m1_coef_rdata[13]),
      .A2F_B_14_3(m1_coef_rdata[12]),
      .A2F_B_14_4(m1_coef_rdata[11]),
      .A2F_B_14_5(m1_coef_rdata[10]),
      .A2F_B_14_6(m1_coef_rdata[9]),
      .A2F_B_14_7(m1_coef_rdata[8]),
      .A2F_B_15_0(m1_coef_rdata[7]),
      .A2F_B_15_1(m1_coef_rdata[6]),
      .A2F_B_15_2(m1_coef_rdata[5]),
      .A2F_B_15_3(m1_coef_rdata[4]),
      .A2F_B_15_4(m1_coef_rdata[3]),
      .A2F_B_15_5(m1_coef_rdata[2]),
      .A2F_B_16_0(m1_coef_rdata[1]),
      .A2F_B_16_1(m1_coef_rdata[0]),
      .A2F_B_16_2(1'b0),
      .A2F_B_16_3(1'b0),
      .A2F_B_16_4(1'b0),
      .A2F_B_16_5(1'b0),
      .A2F_B_16_6(1'b0),
      .A2F_B_16_7(1'b0),
      .A2F_B_17_0(1'b0),
      .A2F_B_17_1(1'b0),
      .A2F_B_17_2(1'b0),
      .A2F_B_17_3(1'b0),
      .A2F_B_17_4(1'b0),
      .A2F_B_17_5(1'b0),
      .A2F_B_18_0(1'b0),
      .A2F_B_18_1(1'b0),
      .A2F_B_18_2(1'b0),
      .A2F_B_18_3(1'b0),
      .A2F_B_18_4(1'b0),
      .A2F_B_18_5(1'b0),
      .A2F_B_18_6(m1_m1_dataout[31]),
      .A2F_B_18_7(m1_m1_dataout[30]),
      .A2F_B_19_0(m1_m1_dataout[29]),
      .A2F_B_19_1(m1_m1_dataout[28]),
      .A2F_B_19_2(m1_m1_dataout[27]),
      .A2F_B_19_3(m1_m1_dataout[26]),
      .A2F_B_19_4(m1_m1_dataout[25]),
      .A2F_B_19_5(m1_m1_dataout[24]),
      .A2F_B_1_0(1'b0),
      .A2F_B_1_1(1'b0),
      .A2F_B_1_2(1'b0),
      .A2F_B_1_3(1'b0),
      .A2F_B_1_4(1'b0),
      .A2F_B_1_5(1'b0),
      .A2F_B_20_0(m1_m1_dataout[23]),
      .A2F_B_20_1(m1_m1_dataout[22]),
      .A2F_B_20_2(m1_m1_dataout[21]),
      .A2F_B_20_3(m1_m1_dataout[20]),
      .A2F_B_20_4(m1_m1_dataout[19]),
      .A2F_B_20_5(m1_m1_dataout[18]),
      .A2F_B_20_6(m1_m1_dataout[17]),
      .A2F_B_20_7(1'b0),
      .A2F_B_21_0(m1_m1_dataout[16]),
      .A2F_B_21_1(m1_m1_dataout[15]),
      .A2F_B_21_2(m1_m1_dataout[14]),
      .A2F_B_21_3(m1_m1_dataout[13]),
      .A2F_B_21_4(m1_m1_dataout[12]),
      .A2F_B_21_5(m1_m1_dataout[11]),
      .A2F_B_22_0(m1_m1_dataout[10]),
      .A2F_B_22_1(m1_m1_dataout[9]),
      .A2F_B_22_2(m1_m1_dataout[8]),
      .A2F_B_22_3(m1_m1_dataout[7]),
      .A2F_B_22_4(m1_m1_dataout[6]),
      .A2F_B_22_5(m1_m1_dataout[5]),
      .A2F_B_22_6(1'b0),
      .A2F_B_22_7(1'b0),
      .A2F_B_23_0(m1_m1_dataout[4]),
      .A2F_B_23_1(m1_m1_dataout[3]),
      .A2F_B_23_2(m1_m1_dataout[2]),
      .A2F_B_23_3(m1_m1_dataout[1]),
      .A2F_B_23_4(m1_m1_dataout[0]),
      .A2F_B_23_5(1'b0),
      .A2F_B_24_0(1'b0),
      .A2F_B_24_1(1'b0),
      .A2F_B_24_2(1'b0),
      .A2F_B_24_3(1'b0),
      .A2F_B_24_4(1'b0),
      .A2F_B_24_5(1'b0),
      .A2F_B_24_6(1'b0),
      .A2F_B_24_7(1'b0),
      .A2F_B_25_0(1'b0),
      .A2F_B_25_1(m1_oper1_rdata[31]),
      .A2F_B_25_2(m1_oper1_rdata[30]),
      .A2F_B_25_3(m1_oper1_rdata[29]),
      .A2F_B_25_4(m1_oper1_rdata[28]),
      .A2F_B_25_5(m1_oper1_rdata[27]),
      .A2F_B_26_0(m1_oper1_rdata[26]),
      .A2F_B_26_1(m1_oper1_rdata[25]),
      .A2F_B_26_2(m1_oper1_rdata[24]),
      .A2F_B_26_3(m1_oper1_rdata[23]),
      .A2F_B_26_4(m1_oper1_rdata[22]),
      .A2F_B_26_5(m1_oper1_rdata[21]),
      .A2F_B_26_6(m1_oper1_rdata[20]),
      .A2F_B_26_7(m1_oper1_rdata[19]),
      .A2F_B_27_0(m1_oper1_rdata[18]),
      .A2F_B_27_1(m1_oper1_rdata[17]),
      .A2F_B_27_2(m1_oper1_rdata[16]),
      .A2F_B_27_3(m1_oper1_rdata[15]),
      .A2F_B_27_4(m1_oper1_rdata[14]),
      .A2F_B_27_5(m1_oper1_rdata[13]),
      .A2F_B_28_0(1'b0),
      .A2F_B_28_1(m1_oper1_rdata[12]),
      .A2F_B_28_2(m1_oper1_rdata[11]),
      .A2F_B_28_3(m1_oper1_rdata[10]),
      .A2F_B_28_4(m1_oper1_rdata[9]),
      .A2F_B_28_5(m1_oper1_rdata[8]),
      .A2F_B_28_6(m1_oper1_rdata[7]),
      .A2F_B_28_7(m1_oper1_rdata[6]),
      .A2F_B_29_0(m1_oper1_rdata[5]),
      .A2F_B_29_1(m1_oper1_rdata[4]),
      .A2F_B_29_2(m1_oper1_rdata[3]),
      .A2F_B_29_3(m1_oper1_rdata[2]),
      .A2F_B_29_4(m1_oper1_rdata[1]),
      .A2F_B_29_5(m1_oper1_rdata[0]),
      .A2F_B_2_0(m1_oper0_rdata[31]),
      .A2F_B_2_1(m1_oper0_rdata[30]),
      .A2F_B_2_2(m1_oper0_rdata[29]),
      .A2F_B_2_3(m1_oper0_rdata[28]),
      .A2F_B_2_4(1'b0),
      .A2F_B_2_5(1'b0),
      .A2F_B_2_6(1'b0),
      .A2F_B_2_7(1'b0),
      .A2F_B_30_0(1'b0),
      .A2F_B_30_1(1'b0),
      .A2F_B_30_2(1'b0),
      .A2F_B_30_3(1'b0),
      .A2F_B_30_4(1'b0),
      .A2F_B_30_5(1'b0),
      .A2F_B_30_6(1'b0),
      .A2F_B_30_7(1'b0),
      .A2F_B_31_0(1'b0),
      .A2F_B_31_1(1'b0),
      .A2F_B_31_2(1'b0),
      .A2F_B_31_3(1'b0),
      .A2F_B_31_4(1'b0),
      .A2F_B_31_5(1'b0),
      .A2F_B_32_0(1'b0),
      .A2F_B_32_1(1'b0),
      .A2F_B_32_2(1'b0),
      .A2F_B_32_3(1'b0),
      .A2F_B_32_4(1'b0),
      .A2F_B_32_5(1'b0),
      .A2F_B_32_6(1'b0),
      .A2F_B_32_7(1'b0),
      .A2F_B_3_0(m1_oper0_rdata[27]),
      .A2F_B_3_1(m1_oper0_rdata[26]),
      .A2F_B_3_2(m1_oper0_rdata[25]),
      .A2F_B_3_3(m1_oper0_rdata[24]),
      .A2F_B_3_4(m1_oper0_rdata[23]),
      .A2F_B_3_5(m1_oper0_rdata[22]),
      .A2F_B_4_0(m1_oper0_rdata[21]),
      .A2F_B_4_1(m1_oper0_rdata[20]),
      .A2F_B_4_2(m1_oper0_rdata[19]),
      .A2F_B_4_3(m1_oper0_rdata[18]),
      .A2F_B_4_4(m1_oper0_rdata[17]),
      .A2F_B_4_5(m1_oper0_rdata[16]),
      .A2F_B_4_6(m1_oper0_rdata[15]),
      .A2F_B_4_7(m1_oper0_rdata[14]),
      .A2F_B_5_0(m1_oper0_rdata[13]),
      .A2F_B_5_1(m1_oper0_rdata[12]),
      .A2F_B_5_2(m1_oper0_rdata[11]),
      .A2F_B_5_3(m1_oper0_rdata[10]),
      .A2F_B_5_4(m1_oper0_rdata[9]),
      .A2F_B_5_5(m1_oper0_rdata[8]),
      .A2F_B_6_0(m1_oper0_rdata[7]),
      .A2F_B_6_1(m1_oper0_rdata[6]),
      .A2F_B_6_2(m1_oper0_rdata[5]),
      .A2F_B_6_3(m1_oper0_rdata[4]),
      .A2F_B_6_4(m1_oper0_rdata[3]),
      .A2F_B_6_5(m1_oper0_rdata[2]),
      .A2F_B_6_6(m1_oper0_rdata[1]),
      .A2F_B_6_7(m1_oper0_rdata[0]),
      .A2F_B_7_0(m1_m0_dataout[31]),
      .A2F_B_7_1(m1_m0_dataout[30]),
      .A2F_B_7_2(m1_m0_dataout[29]),
      .A2F_B_7_3(m1_m0_dataout[28]),
      .A2F_B_7_4(m1_m0_dataout[27]),
      .A2F_B_7_5(m1_m0_dataout[26]),
      .A2F_B_8_0(m1_m0_dataout[25]),
      .A2F_B_8_1(m1_m0_dataout[24]),
      .A2F_B_8_2(m1_m0_dataout[23]),
      .A2F_B_8_3(m1_m0_dataout[22]),
      .A2F_B_8_4(m1_m0_dataout[21]),
      .A2F_B_8_5(m1_m0_dataout[20]),
      .A2F_B_8_6(m1_m0_dataout[19]),
      .A2F_B_8_7(m1_m0_dataout[18]),
      .A2F_B_9_0(m1_m0_dataout[17]),
      .A2F_B_9_1(m1_m0_dataout[16]),
      .A2F_B_9_2(m1_m0_dataout[15]),
      .A2F_B_9_3(m1_m0_dataout[14]),
      .A2F_B_9_4(m1_m0_dataout[13]),
      .A2F_B_9_5(m1_m0_dataout[12]),
      .A2F_L_10_0(lint_WDATA[16]),
      .A2F_L_10_1(lint_WDATA[17]),
      .A2F_L_10_2(lint_WDATA[18]),
      .A2F_L_10_3(lint_WDATA[19]),
      .A2F_L_10_4(lint_WDATA[20]),
      .A2F_L_10_5(lint_WDATA[21]),
      .A2F_L_10_6(lint_WDATA[22]),
      .A2F_L_10_7(lint_WDATA[23]),
      .A2F_L_11_0(lint_WDATA[24]),
      .A2F_L_11_1(lint_WDATA[25]),
      .A2F_L_11_2(lint_WDATA[26]),
      .A2F_L_11_3(lint_WDATA[27]),
      .A2F_L_11_4(lint_WDATA[28]),
      .A2F_L_11_5(lint_WDATA[29]),
      .A2F_L_12_0(lint_WDATA[30]),
      .A2F_L_12_1(lint_WDATA[31]),
      .A2F_L_12_2(lint_REQ),
      .A2F_L_12_3(lint_WEN),
      .A2F_L_12_4(lint_BE[0]),
      .A2F_L_12_5(lint_BE[1]),
      .A2F_L_12_6(lint_BE[2]),
      .A2F_L_12_7(lint_BE[3]),
      .A2F_L_13_0(lint_ADDR[0]),
      .A2F_L_13_1(lint_ADDR[1]),
      .A2F_L_13_2(lint_ADDR[2]),
      .A2F_L_13_3(lint_ADDR[3]),
      .A2F_L_13_4(lint_ADDR[4]),
      .A2F_L_13_5(lint_ADDR[5]),
      .A2F_L_14_0(lint_ADDR[6]),
      .A2F_L_14_1(lint_ADDR[7]),
      .A2F_L_14_2(lint_ADDR[8]),
      .A2F_L_14_3(lint_ADDR[9]),
      .A2F_L_14_4(lint_ADDR[10]),
      .A2F_L_14_5(lint_ADDR[11]),
      .A2F_L_14_6(lint_ADDR[12]),
      .A2F_L_14_7(lint_ADDR[13]),
      .A2F_L_15_0(lint_ADDR[14]),
      .A2F_L_15_1(lint_ADDR[15]),
      .A2F_L_15_2(lint_ADDR[16]),
      .A2F_L_15_3(lint_ADDR[17]),
      .A2F_L_15_4(lint_ADDR[18]),
      .A2F_L_15_5(lint_ADDR[19]),
      .A2F_L_16_0(fpgaio_in[64]),
      .A2F_L_16_1(fpgaio_in[65]),
      .A2F_L_16_2(fpgaio_in[66]),
      .A2F_L_16_3(fpgaio_in[67]),
      .A2F_L_16_4(fpgaio_in[68]),
      .A2F_L_16_5(fpgaio_in[69]),
      .A2F_L_16_6(fpgaio_in[70]),
      .A2F_L_16_7(fpgaio_in[71]),
      .A2F_L_17_0(fpgaio_in[72]),
      .A2F_L_17_1(fpgaio_in[73]),
      .A2F_L_17_2(fpgaio_in[74]),
      .A2F_L_17_3(fpgaio_in[75]),
      .A2F_L_17_4(fpgaio_in[76]),
      .A2F_L_17_5(fpgaio_in[77]),
      .A2F_L_18_0(fpgaio_in[78]),
      .A2F_L_18_1(fpgaio_in[79]),
      .A2F_L_18_2(1'b0),
      .A2F_L_18_3(1'b0),
      .A2F_L_18_4(1'b0),
      .A2F_L_18_5(1'b0),
      .A2F_L_18_6(1'b0),
      .A2F_L_18_7(1'b0),
      .A2F_L_19_0(control_in[0]),
      .A2F_L_19_1(control_in[1]),
      .A2F_L_19_2(control_in[2]),
      .A2F_L_19_3(control_in[3]),
      .A2F_L_19_4(control_in[4]),
      .A2F_L_19_5(control_in[5]),
      .A2F_L_1_0(1'b0),
      .A2F_L_1_1(1'b0),
      .A2F_L_1_2(1'b0),
      .A2F_L_1_3(1'b0),
      .A2F_L_1_4(1'b0),
      .A2F_L_1_5(1'b0),
      .A2F_L_20_0(control_in[6]),
      .A2F_L_20_1(control_in[7]),
      .A2F_L_20_2(control_in[8]),
      .A2F_L_20_3(control_in[9]),
      .A2F_L_20_4(control_in[10]),
      .A2F_L_20_5(control_in[11]),
      .A2F_L_20_6(control_in[12]),
      .A2F_L_20_7(control_in[13]),
      .A2F_L_21_0(control_in[14]),
      .A2F_L_21_1(control_in[15]),
      .A2F_L_21_2(control_in[16]),
      .A2F_L_21_3(control_in[17]),
      .A2F_L_21_4(control_in[18]),
      .A2F_L_21_5(control_in[19]),
      .A2F_L_22_0(control_in[20]),
      .A2F_L_22_1(control_in[21]),
      .A2F_L_22_2(control_in[22]),
      .A2F_L_22_3(control_in[23]),
      .A2F_L_22_4(control_in[24]),
      .A2F_L_22_5(control_in[25]),
      .A2F_L_22_6(control_in[26]),
      .A2F_L_22_7(1'b0),
      .A2F_L_23_0(control_in[27]),
      .A2F_L_23_1(control_in[28]),
      .A2F_L_23_2(control_in[29]),
      .A2F_L_23_3(control_in[30]),
      .A2F_L_23_4(control_in[31]),
      .A2F_L_23_5(1'b0),
      .A2F_L_24_0(1'b0),
      .A2F_L_24_1(1'b0),
      .A2F_L_24_2(1'b0),
      .A2F_L_24_3(1'b0),
      .A2F_L_24_4(1'b0),
      .A2F_L_24_5(1'b0),
      .A2F_L_24_6(1'b0),
      .A2F_L_24_7(1'b0),
      .A2F_L_25_0(fpgaio_in[32]),
      .A2F_L_25_1(fpgaio_in[33]),
      .A2F_L_25_2(RESET[3]),
      .A2F_L_25_3(fpgaio_in[34]),
      .A2F_L_25_4(fpgaio_in[35]),
      .A2F_L_25_5(1'b0),
      .A2F_L_26_0(fpgaio_in[36]),
      .A2F_L_26_1(fpgaio_in[37]),
      .A2F_L_26_2(fpgaio_in[38]),
      .A2F_L_26_3(fpgaio_in[39]),
      .A2F_L_26_4(1'b0),
      .A2F_L_26_5(1'b0),
      .A2F_L_26_6(1'b0),
      .A2F_L_26_7(1'b0),
      .A2F_L_27_0(fpgaio_in[40]),
      .A2F_L_27_1(fpgaio_in[41]),
      .A2F_L_27_2(fpgaio_in[42]),
      .A2F_L_27_3(fpgaio_in[43]),
      .A2F_L_27_4(1'b0),
      .A2F_L_27_5(1'b0),
      .A2F_L_28_0(fpgaio_in[44]),
      .A2F_L_28_1(fpgaio_in[45]),
      .A2F_L_28_2(fpgaio_in[46]),
      .A2F_L_28_3(fpgaio_in[47]),
      .A2F_L_28_4(1'b0),
      .A2F_L_28_5(1'b0),
      .A2F_L_28_6(1'b0),
      .A2F_L_28_7(1'b0),
      .A2F_L_29_0(fpgaio_in[48]),
      .A2F_L_29_1(fpgaio_in[49]),
      .A2F_L_29_2(fpgaio_in[50]),
      .A2F_L_29_3(fpgaio_in[51]),
      .A2F_L_29_4(1'b0),
      .A2F_L_29_5(1'b0),
      .A2F_L_2_0(fpgaio_in[0]),
      .A2F_L_2_1(fpgaio_in[1]),
      .A2F_L_2_2(fpgaio_in[2]),
      .A2F_L_2_3(fpgaio_in[3]),
      .A2F_L_2_4(RESET[0]),
      .A2F_L_2_5(1'b0),
      .A2F_L_2_6(1'b0),
      .A2F_L_2_7(1'b0),
      .A2F_L_30_0(fpgaio_in[52]),
      .A2F_L_30_1(fpgaio_in[53]),
      .A2F_L_30_2(fpgaio_in[54]),
      .A2F_L_30_3(fpgaio_in[55]),
      .A2F_L_30_4(1'b0),
      .A2F_L_30_5(1'b0),
      .A2F_L_30_6(1'b0),
      .A2F_L_30_7(1'b0),
      .A2F_L_31_0(fpgaio_in[56]),
      .A2F_L_31_1(fpgaio_in[57]),
      .A2F_L_31_2(fpgaio_in[58]),
      .A2F_L_31_3(fpgaio_in[59]),
      .A2F_L_31_4(1'b0),
      .A2F_L_31_5(1'b0),
      .A2F_L_32_0(fpgaio_in[60]),
      .A2F_L_32_1(fpgaio_in[61]),
      .A2F_L_32_2(fpgaio_in[62]),
      .A2F_L_32_3(fpgaio_in[63]),
      .A2F_L_32_4(1'b0),
      .A2F_L_32_5(1'b0),
      .A2F_L_32_6(1'b0),
      .A2F_L_32_7(1'b0),
      .A2F_L_3_0(fpgaio_in[4]),
      .A2F_L_3_1(fpgaio_in[5]),
      .A2F_L_3_2(fpgaio_in[6]),
      .A2F_L_3_3(fpgaio_in[7]),
      .A2F_L_3_4(fpgaio_in[8]),
      .A2F_L_3_5(fpgaio_in[9]),
      .A2F_L_4_0(1'b0),
      .A2F_L_4_1(1'b0),
      .A2F_L_4_2(fpgaio_in[10]),
      .A2F_L_4_3(fpgaio_in[11]),
      .A2F_L_4_4(fpgaio_in[12]),
      .A2F_L_4_5(fpgaio_in[13]),
      .A2F_L_4_6(fpgaio_in[14]),
      .A2F_L_4_7(fpgaio_in[15]),
      .A2F_L_5_0(fpgaio_in[16]),
      .A2F_L_5_1(fpgaio_in[17]),
      .A2F_L_5_2(fpgaio_in[18]),
      .A2F_L_5_3(fpgaio_in[19]),
      .A2F_L_5_4(fpgaio_in[20]),
      .A2F_L_5_5(fpgaio_in[21]),
      .A2F_L_6_0(fpgaio_in[22]),
      .A2F_L_6_1(fpgaio_in[23]),
      .A2F_L_6_2(fpgaio_in[24]),
      .A2F_L_6_3(fpgaio_in[25]),
      .A2F_L_6_4(fpgaio_in[26]),
      .A2F_L_6_5(fpgaio_in[27]),
      .A2F_L_6_6(1'b0),
      .A2F_L_6_7(1'b0),
      .A2F_L_7_0(fpgaio_in[28]),
      .A2F_L_7_1(fpgaio_in[29]),
      .A2F_L_7_2(fpgaio_in[30]),
      .A2F_L_7_3(fpgaio_in[31]),
      .A2F_L_7_4(lint_WDATA[0]),
      .A2F_L_7_5(lint_WDATA[1]),
      .A2F_L_8_0(lint_WDATA[2]),
      .A2F_L_8_1(lint_WDATA[3]),
      .A2F_L_8_2(lint_WDATA[4]),
      .A2F_L_8_3(lint_WDATA[5]),
      .A2F_L_8_4(lint_WDATA[6]),
      .A2F_L_8_5(lint_WDATA[7]),
      .A2F_L_8_6(lint_WDATA[8]),
      .A2F_L_8_7(lint_WDATA[9]),
      .A2F_L_9_0(lint_WDATA[10]),
      .A2F_L_9_1(lint_WDATA[11]),
      .A2F_L_9_2(lint_WDATA[12]),
      .A2F_L_9_3(lint_WDATA[13]),
      .A2F_L_9_4(lint_WDATA[14]),
      .A2F_L_9_5(lint_WDATA[15]),
      .A2F_T_10_0(tcdm_rdata_p1[4]),
      .A2F_T_10_1(tcdm_rdata_p1[5]),
      .A2F_T_10_2(tcdm_rdata_p1[6]),
      .A2F_T_10_3(tcdm_rdata_p1[7]),
      .A2F_T_10_4(tcdm_rdata_p1[8]),
      .A2F_T_10_5(tcdm_rdata_p1[9]),
      .A2F_T_10_6(tcdm_rdata_p1[10]),
      .A2F_T_10_7(tcdm_rdata_p1[11]),
      .A2F_T_11_0(tcdm_rdata_p1[12]),
      .A2F_T_11_1(tcdm_rdata_p1[13]),
      .A2F_T_11_2(tcdm_rdata_p1[14]),
      .A2F_T_11_3(tcdm_rdata_p1[15]),
      .A2F_T_11_4(tcdm_fmo_p1),
      .A2F_T_11_5(1'b0),
      .A2F_T_12_0(1'b0),
      .A2F_T_12_1(tcdm_rdata_p1[16]),
      .A2F_T_12_2(tcdm_rdata_p1[17]),
      .A2F_T_12_3(tcdm_rdata_p1[18]),
      .A2F_T_12_4(tcdm_rdata_p1[19]),
      .A2F_T_12_5(tcdm_rdata_p1[20]),
      .A2F_T_12_6(tcdm_rdata_p1[21]),
      .A2F_T_12_7(1'b0),
      .A2F_T_13_0(tcdm_rdata_p1[22]),
      .A2F_T_13_1(tcdm_rdata_p1[23]),
      .A2F_T_13_2(tcdm_rdata_p1[24]),
      .A2F_T_13_3(tcdm_rdata_p1[25]),
      .A2F_T_13_4(tcdm_rdata_p1[26]),
      .A2F_T_13_5(tcdm_rdata_p1[27]),
      .A2F_T_14_0(tcdm_rdata_p1[28]),
      .A2F_T_14_1(tcdm_rdata_p1[29]),
      .A2F_T_14_2(tcdm_rdata_p1[30]),
      .A2F_T_14_3(tcdm_rdata_p1[31]),
      .A2F_T_14_4(1'b0),
      .A2F_T_14_5(1'b0),
      .A2F_T_14_6(1'b0),
      .A2F_T_14_7(1'b0),
      .A2F_T_15_0(1'b0),
      .A2F_T_15_1(1'b0),
      .A2F_T_15_2(1'b0),
      .A2F_T_15_3(1'b0),
      .A2F_T_15_4(1'b0),
      .A2F_T_15_5(1'b0),
      .A2F_T_16_0(1'b0),
      .A2F_T_16_1(1'b0),
      .A2F_T_16_2(1'b0),
      .A2F_T_16_3(1'b0),
      .A2F_T_16_4(1'b0),
      .A2F_T_16_5(1'b0),
      .A2F_T_16_6(1'b0),
      .A2F_T_16_7(1'b0),
      .A2F_T_17_0(tcdm_rdata_p2[0]),
      .A2F_T_17_1(tcdm_rdata_p2[1]),
      .A2F_T_17_2(tcdm_rdata_p2[2]),
      .A2F_T_17_3(tcdm_rdata_p2[3]),
      .A2F_T_17_4(tcdm_valid_p2),
      .A2F_T_17_5(tcdm_gnt_p2),
      .A2F_T_18_0(tcdm_rdata_p2[4]),
      .A2F_T_18_1(tcdm_rdata_p2[5]),
      .A2F_T_18_2(tcdm_rdata_p2[6]),
      .A2F_T_18_3(tcdm_rdata_p2[7]),
      .A2F_T_18_4(tcdm_rdata_p2[8]),
      .A2F_T_18_5(tcdm_rdata_p2[9]),
      .A2F_T_18_6(tcdm_rdata_p2[10]),
      .A2F_T_18_7(tcdm_rdata_p2[11]),
      .A2F_T_19_0(tcdm_rdata_p2[12]),
      .A2F_T_19_1(tcdm_rdata_p2[13]),
      .A2F_T_19_2(tcdm_rdata_p2[14]),
      .A2F_T_19_3(tcdm_rdata_p2[15]),
      .A2F_T_19_4(tcdm_fmo_p2),
      .A2F_T_19_5(1'b0),
      .A2F_T_1_0(1'b0),
      .A2F_T_1_1(1'b0),
      .A2F_T_1_2(1'b0),
      .A2F_T_1_3(1'b0),
      .A2F_T_1_4(1'b0),
      .A2F_T_1_5(1'b0),
      .A2F_T_20_0(1'b0),
      .A2F_T_20_1(tcdm_rdata_p2[16]),
      .A2F_T_20_2(tcdm_rdata_p2[17]),
      .A2F_T_20_3(tcdm_rdata_p2[18]),
      .A2F_T_20_4(tcdm_rdata_p2[19]),
      .A2F_T_20_5(tcdm_rdata_p2[20]),
      .A2F_T_20_6(tcdm_rdata_p2[21]),
      .A2F_T_20_7(1'b0),
      .A2F_T_21_0(tcdm_rdata_p2[22]),
      .A2F_T_21_1(tcdm_rdata_p2[23]),
      .A2F_T_21_2(tcdm_rdata_p2[24]),
      .A2F_T_21_3(tcdm_rdata_p2[25]),
      .A2F_T_21_4(tcdm_rdata_p2[26]),
      .A2F_T_21_5(tcdm_rdata_p2[27]),
      .A2F_T_22_0(tcdm_rdata_p2[28]),
      .A2F_T_22_1(tcdm_rdata_p2[29]),
      .A2F_T_22_2(tcdm_rdata_p2[30]),
      .A2F_T_22_3(tcdm_rdata_p2[31]),
      .A2F_T_22_4(1'b0),
      .A2F_T_22_5(1'b0),
      .A2F_T_22_6(1'b0),
      .A2F_T_22_7(1'b0),
      .A2F_T_23_0(tcdm_rdata_p3[0]),
      .A2F_T_23_1(tcdm_rdata_p3[1]),
      .A2F_T_23_2(tcdm_rdata_p3[2]),
      .A2F_T_23_3(tcdm_rdata_p3[3]),
      .A2F_T_23_4(tcdm_valid_p3),
      .A2F_T_23_5(tcdm_gnt_p3),
      .A2F_T_24_0(tcdm_rdata_p3[4]),
      .A2F_T_24_1(tcdm_rdata_p3[5]),
      .A2F_T_24_2(tcdm_rdata_p3[6]),
      .A2F_T_24_3(tcdm_rdata_p3[7]),
      .A2F_T_24_4(tcdm_rdata_p3[8]),
      .A2F_T_24_5(tcdm_rdata_p3[9]),
      .A2F_T_24_6(tcdm_rdata_p3[10]),
      .A2F_T_24_7(tcdm_rdata_p3[11]),
      .A2F_T_25_0(tcdm_rdata_p3[12]),
      .A2F_T_25_1(tcdm_rdata_p3[13]),
      .A2F_T_25_2(tcdm_rdata_p3[14]),
      .A2F_T_25_3(tcdm_rdata_p3[15]),
      .A2F_T_25_4(tcdm_fmo_p3),
      .A2F_T_25_5(1'b0),
      .A2F_T_26_0(1'b0),
      .A2F_T_26_1(tcdm_rdata_p3[16]),
      .A2F_T_26_2(tcdm_rdata_p3[17]),
      .A2F_T_26_3(tcdm_rdata_p3[18]),
      .A2F_T_26_4(tcdm_rdata_p3[19]),
      .A2F_T_26_5(tcdm_rdata_p3[20]),
      .A2F_T_26_6(tcdm_rdata_p3[21]),
      .A2F_T_26_7(1'b0),
      .A2F_T_27_0(tcdm_rdata_p3[22]),
      .A2F_T_27_1(tcdm_rdata_p3[23]),
      .A2F_T_27_2(tcdm_rdata_p3[24]),
      .A2F_T_27_3(tcdm_rdata_p3[25]),
      .A2F_T_27_4(tcdm_rdata_p3[26]),
      .A2F_T_27_5(tcdm_rdata_p3[27]),
      .A2F_T_28_0(tcdm_rdata_p3[28]),
      .A2F_T_28_1(tcdm_rdata_p3[29]),
      .A2F_T_28_2(tcdm_rdata_p3[30]),
      .A2F_T_28_3(tcdm_rdata_p3[31]),
      .A2F_T_28_4(1'b0),
      .A2F_T_28_5(1'b0),
      .A2F_T_28_6(1'b0),
      .A2F_T_28_7(1'b0),
      .A2F_T_29_0(1'b0),
      .A2F_T_29_1(1'b0),
      .A2F_T_29_2(RESET[2]),
      .A2F_T_29_3(1'b0),
      .A2F_T_29_4(1'b0),
      .A2F_T_29_5(1'b0),
      .A2F_T_2_0(1'b0),
      .A2F_T_2_1(1'b0),
      .A2F_T_2_2(1'b0),
      .A2F_T_2_3(1'b0),
      .A2F_T_2_4(1'b0),
      .A2F_T_2_5(1'b0),
      .A2F_T_2_6(1'b0),
      .A2F_T_2_7(1'b0),
      .A2F_T_30_0(1'b0),
      .A2F_T_30_1(1'b0),
      .A2F_T_30_2(1'b0),
      .A2F_T_30_3(1'b0),
      .A2F_T_30_4(1'b0),
      .A2F_T_30_5(1'b0),
      .A2F_T_30_6(1'b0),
      .A2F_T_30_7(1'b0),
      .A2F_T_31_0(1'b0),
      .A2F_T_31_1(1'b0),
      .A2F_T_31_2(1'b0),
      .A2F_T_31_3(1'b0),
      .A2F_T_31_4(1'b0),
      .A2F_T_31_5(1'b0),
      .A2F_T_32_0(1'b0),
      .A2F_T_32_1(1'b0),
      .A2F_T_32_2(1'b0),
      .A2F_T_32_3(1'b0),
      .A2F_T_32_4(1'b0),
      .A2F_T_32_5(1'b0),
      .A2F_T_32_6(1'b0),
      .A2F_T_32_7(1'b0),
      .A2F_T_3_0(tcdm_rdata_p0[0]),
      .A2F_T_3_1(tcdm_rdata_p0[1]),
      .A2F_T_3_2(tcdm_rdata_p0[2]),
      .A2F_T_3_3(tcdm_rdata_p0[3]),
      .A2F_T_3_4(tcdm_valid_p0),
      .A2F_T_3_5(tcdm_gnt_p0),
      .A2F_T_4_0(tcdm_rdata_p0[4]),
      .A2F_T_4_1(tcdm_rdata_p0[5]),
      .A2F_T_4_2(tcdm_rdata_p0[6]),
      .A2F_T_4_3(tcdm_rdata_p0[7]),
      .A2F_T_4_4(tcdm_rdata_p0[8]),
      .A2F_T_4_5(tcdm_rdata_p0[9]),
      .A2F_T_4_6(tcdm_rdata_p0[10]),
      .A2F_T_4_7(tcdm_rdata_p0[11]),
      .A2F_T_5_0(tcdm_rdata_p0[12]),
      .A2F_T_5_1(tcdm_rdata_p0[13]),
      .A2F_T_5_2(tcdm_rdata_p0[14]),
      .A2F_T_5_3(tcdm_rdata_p0[15]),
      .A2F_T_5_4(tcdm_fmo_p0),
      .A2F_T_5_5(1'b0),
      .A2F_T_6_0(RESET[1]),
      .A2F_T_6_1(tcdm_rdata_p0[16]),
      .A2F_T_6_2(tcdm_rdata_p0[17]),
      .A2F_T_6_3(tcdm_rdata_p0[18]),
      .A2F_T_6_4(tcdm_rdata_p0[19]),
      .A2F_T_6_5(tcdm_rdata_p0[20]),
      .A2F_T_6_6(tcdm_rdata_p0[21]),
      .A2F_T_6_7(1'b0),
      .A2F_T_7_0(tcdm_rdata_p0[22]),
      .A2F_T_7_1(tcdm_rdata_p0[23]),
      .A2F_T_7_2(tcdm_rdata_p0[24]),
      .A2F_T_7_3(tcdm_rdata_p0[25]),
      .A2F_T_7_4(tcdm_rdata_p0[26]),
      .A2F_T_7_5(tcdm_rdata_p0[27]),
      .A2F_T_8_0(tcdm_rdata_p0[28]),
      .A2F_T_8_1(tcdm_rdata_p0[29]),
      .A2F_T_8_2(tcdm_rdata_p0[30]),
      .A2F_T_8_3(tcdm_rdata_p0[31]),
      .A2F_T_8_4(1'b0),
      .A2F_T_8_5(1'b0),
      .A2F_T_8_6(1'b0),
      .A2F_T_8_7(1'b0),
      .A2F_T_9_0(tcdm_rdata_p1[0]),
      .A2F_T_9_1(tcdm_rdata_p1[1]),
      .A2F_T_9_2(tcdm_rdata_p1[2]),
      .A2F_T_9_3(tcdm_rdata_p1[3]),
      .A2F_T_9_4(tcdm_valid_p1),
      .A2F_T_9_5(tcdm_gnt_p1),
      .A2F_R_10_0(m0_m0_dataout[11]),
      .A2F_R_10_1(m0_m0_dataout[10]),
      .A2F_R_10_2(m0_m0_dataout[9]),
      .A2F_R_10_3(m0_m0_dataout[8]),
      .A2F_R_10_4(m0_m0_dataout[7]),
      .A2F_R_10_5(m0_m0_dataout[6]),
      .A2F_R_10_6(m0_m0_dataout[5]),
      .A2F_R_10_7(m0_m0_dataout[4]),
      .A2F_R_11_0(m0_m0_dataout[3]),
      .A2F_R_11_1(m0_m0_dataout[2]),
      .A2F_R_11_2(m0_m0_dataout[1]),
      .A2F_R_11_3(m0_m0_dataout[0]),
      .A2F_R_11_4(m0_coef_rdata[31]),
      .A2F_R_11_5(m0_coef_rdata[30]),
      .A2F_R_12_0(m0_coef_rdata[29]),
      .A2F_R_12_1(m0_coef_rdata[28]),
      .A2F_R_12_2(m0_coef_rdata[27]),
      .A2F_R_12_3(m0_coef_rdata[26]),
      .A2F_R_12_4(m0_coef_rdata[25]),
      .A2F_R_12_5(m0_coef_rdata[24]),
      .A2F_R_12_6(m0_coef_rdata[23]),
      .A2F_R_12_7(m0_coef_rdata[22]),
      .A2F_R_13_0(m0_coef_rdata[21]),
      .A2F_R_13_1(m0_coef_rdata[20]),
      .A2F_R_13_2(m0_coef_rdata[19]),
      .A2F_R_13_3(m0_coef_rdata[18]),
      .A2F_R_13_4(m0_coef_rdata[17]),
      .A2F_R_13_5(m0_coef_rdata[16]),
      .A2F_R_14_0(m0_coef_rdata[15]),
      .A2F_R_14_1(m0_coef_rdata[14]),
      .A2F_R_14_2(m0_coef_rdata[13]),
      .A2F_R_14_3(m0_coef_rdata[12]),
      .A2F_R_14_4(m0_coef_rdata[11]),
      .A2F_R_14_5(m0_coef_rdata[10]),
      .A2F_R_14_6(m0_coef_rdata[9]),
      .A2F_R_14_7(m0_coef_rdata[8]),
      .A2F_R_15_0(m0_coef_rdata[7]),
      .A2F_R_15_1(m0_coef_rdata[6]),
      .A2F_R_15_2(m0_coef_rdata[5]),
      .A2F_R_15_3(m0_coef_rdata[4]),
      .A2F_R_15_4(m0_coef_rdata[3]),
      .A2F_R_15_5(m0_coef_rdata[2]),
      .A2F_R_16_0(m0_coef_rdata[1]),
      .A2F_R_16_1(m0_coef_rdata[0]),
      .A2F_R_16_2(1'b0),
      .A2F_R_16_3(1'b0),
      .A2F_R_16_4(1'b0),
      .A2F_R_16_5(1'b0),
      .A2F_R_16_6(1'b0),
      .A2F_R_16_7(1'b0),
      .A2F_R_17_0(1'b0),
      .A2F_R_17_1(1'b0),
      .A2F_R_17_2(1'b0),
      .A2F_R_17_3(1'b0),
      .A2F_R_17_4(1'b0),
      .A2F_R_17_5(1'b0),
      .A2F_R_18_0(m0_m1_dataout[31]),
      .A2F_R_18_1(m0_m1_dataout[30]),
      .A2F_R_18_2(m0_m1_dataout[29]),
      .A2F_R_18_3(m0_m1_dataout[28]),
      .A2F_R_18_4(m0_m1_dataout[27]),
      .A2F_R_18_5(m0_m1_dataout[26]),
      .A2F_R_18_6(m0_m1_dataout[25]),
      .A2F_R_18_7(m0_m1_dataout[24]),
      .A2F_R_19_0(m0_m1_dataout[23]),
      .A2F_R_19_1(m0_m1_dataout[22]),
      .A2F_R_19_2(m0_m1_dataout[21]),
      .A2F_R_19_3(m0_m1_dataout[20]),
      .A2F_R_19_4(m0_m1_dataout[19]),
      .A2F_R_19_5(m0_m1_dataout[18]),
      .A2F_R_1_0(1'b0),
      .A2F_R_1_1(1'b0),
      .A2F_R_1_2(1'b0),
      .A2F_R_1_3(1'b0),
      .A2F_R_1_4(1'b0),
      .A2F_R_1_5(1'b0),
      .A2F_R_20_0(m0_m1_dataout[17]),
      .A2F_R_20_1(m0_m1_dataout[16]),
      .A2F_R_20_2(m0_m1_dataout[15]),
      .A2F_R_20_3(m0_m1_dataout[14]),
      .A2F_R_20_4(m0_m1_dataout[13]),
      .A2F_R_20_5(m0_m1_dataout[12]),
      .A2F_R_20_6(m0_m1_dataout[11]),
      .A2F_R_20_7(1'b0),
      .A2F_R_21_0(m0_m1_dataout[10]),
      .A2F_R_21_1(m0_m1_dataout[9]),
      .A2F_R_21_2(m0_m1_dataout[8]),
      .A2F_R_21_3(m0_m1_dataout[7]),
      .A2F_R_21_4(m0_m1_dataout[6]),
      .A2F_R_21_5(m0_m1_dataout[5]),
      .A2F_R_22_0(m0_m1_dataout[4]),
      .A2F_R_22_1(m0_m1_dataout[3]),
      .A2F_R_22_2(m0_m1_dataout[2]),
      .A2F_R_22_3(m0_m1_dataout[1]),
      .A2F_R_22_4(m0_m1_dataout[0]),
      .A2F_R_22_5(1'b0),
      .A2F_R_22_6(1'b0),
      .A2F_R_22_7(1'b0),
      .A2F_R_23_0(1'b0),
      .A2F_R_23_1(1'b0),
      .A2F_R_23_2(1'b0),
      .A2F_R_23_3(1'b0),
      .A2F_R_23_4(1'b0),
      .A2F_R_23_5(1'b0),
      .A2F_R_24_0(1'b0),
      .A2F_R_24_1(1'b0),
      .A2F_R_24_2(1'b0),
      .A2F_R_24_3(1'b0),
      .A2F_R_24_4(1'b0),
      .A2F_R_24_5(1'b0),
      .A2F_R_24_6(1'b0),
      .A2F_R_24_7(1'b0),
      .A2F_R_25_0(1'b0),
      .A2F_R_25_1(m0_oper1_rdata[31]),
      .A2F_R_25_2(m0_oper1_rdata[30]),
      .A2F_R_25_3(m0_oper1_rdata[29]),
      .A2F_R_25_4(m0_oper1_rdata[28]),
      .A2F_R_25_5(m0_oper1_rdata[27]),
      .A2F_R_26_0(m0_oper1_rdata[26]),
      .A2F_R_26_1(m0_oper1_rdata[25]),
      .A2F_R_26_2(m0_oper1_rdata[24]),
      .A2F_R_26_3(m0_oper1_rdata[23]),
      .A2F_R_26_4(m0_oper1_rdata[22]),
      .A2F_R_26_5(m0_oper1_rdata[21]),
      .A2F_R_26_6(m0_oper1_rdata[20]),
      .A2F_R_26_7(m0_oper1_rdata[19]),
      .A2F_R_27_0(m0_oper1_rdata[18]),
      .A2F_R_27_1(m0_oper1_rdata[17]),
      .A2F_R_27_2(m0_oper1_rdata[16]),
      .A2F_R_27_3(m0_oper1_rdata[15]),
      .A2F_R_27_4(m0_oper1_rdata[14]),
      .A2F_R_27_5(m0_oper1_rdata[13]),
      .A2F_R_28_0(1'b0),
      .A2F_R_28_1(m0_oper1_rdata[12]),
      .A2F_R_28_2(m0_oper1_rdata[11]),
      .A2F_R_28_3(m0_oper1_rdata[10]),
      .A2F_R_28_4(m0_oper1_rdata[9]),
      .A2F_R_28_5(m0_oper1_rdata[8]),
      .A2F_R_28_6(m0_oper1_rdata[7]),
      .A2F_R_28_7(m0_oper1_rdata[6]),
      .A2F_R_29_0(m0_oper1_rdata[5]),
      .A2F_R_29_1(m0_oper1_rdata[4]),
      .A2F_R_29_2(m0_oper1_rdata[3]),
      .A2F_R_29_3(m0_oper1_rdata[2]),
      .A2F_R_29_4(m0_oper1_rdata[1]),
      .A2F_R_29_5(m0_oper1_rdata[0]),
      .A2F_R_2_0(m0_oper0_rdata[31]),
      .A2F_R_2_1(m0_oper0_rdata[30]),
      .A2F_R_2_2(m0_oper0_rdata[29]),
      .A2F_R_2_3(m0_oper0_rdata[28]),
      .A2F_R_2_4(1'b0),
      .A2F_R_2_5(1'b0),
      .A2F_R_2_6(1'b0),
      .A2F_R_2_7(1'b0),
      .A2F_R_30_0(1'b0),
      .A2F_R_30_1(1'b0),
      .A2F_R_30_2(1'b0),
      .A2F_R_30_3(1'b0),
      .A2F_R_30_4(1'b0),
      .A2F_R_30_5(1'b0),
      .A2F_R_30_6(1'b0),
      .A2F_R_30_7(1'b0),
      .A2F_R_31_0(1'b0),
      .A2F_R_31_1(1'b0),
      .A2F_R_31_2(1'b0),
      .A2F_R_31_3(1'b0),
      .A2F_R_31_4(1'b0),
      .A2F_R_31_5(1'b0),
      .A2F_R_32_0(1'b0),
      .A2F_R_32_1(1'b0),
      .A2F_R_32_2(1'b0),
      .A2F_R_32_3(1'b0),
      .A2F_R_32_4(1'b0),
      .A2F_R_32_5(1'b0),
      .A2F_R_32_6(1'b0),
      .A2F_R_32_7(1'b0),
      .A2F_R_3_0(m0_oper0_rdata[27]),
      .A2F_R_3_1(m0_oper0_rdata[26]),
      .A2F_R_3_2(m0_oper0_rdata[25]),
      .A2F_R_3_3(m0_oper0_rdata[24]),
      .A2F_R_3_4(m0_oper0_rdata[23]),
      .A2F_R_3_5(m0_oper0_rdata[22]),
      .A2F_R_4_0(m0_oper0_rdata[21]),
      .A2F_R_4_1(m0_oper0_rdata[20]),
      .A2F_R_4_2(m0_oper0_rdata[19]),
      .A2F_R_4_3(m0_oper0_rdata[18]),
      .A2F_R_4_4(m0_oper0_rdata[17]),
      .A2F_R_4_5(m0_oper0_rdata[16]),
      .A2F_R_4_6(m0_oper0_rdata[15]),
      .A2F_R_4_7(m0_oper0_rdata[14]),
      .A2F_R_5_0(m0_oper0_rdata[13]),
      .A2F_R_5_1(m0_oper0_rdata[12]),
      .A2F_R_5_2(m0_oper0_rdata[11]),
      .A2F_R_5_3(m0_oper0_rdata[10]),
      .A2F_R_5_4(m0_oper0_rdata[9]),
      .A2F_R_5_5(m0_oper0_rdata[8]),
      .A2F_R_6_0(m0_oper0_rdata[7]),
      .A2F_R_6_1(m0_oper0_rdata[6]),
      .A2F_R_6_2(m0_oper0_rdata[5]),
      .A2F_R_6_3(m0_oper0_rdata[4]),
      .A2F_R_6_4(m0_oper0_rdata[3]),
      .A2F_R_6_5(m0_oper0_rdata[2]),
      .A2F_R_6_6(m0_oper0_rdata[1]),
      .A2F_R_6_7(m0_oper0_rdata[0]),
      .A2F_R_7_0(m0_m0_dataout[31]),
      .A2F_R_7_1(m0_m0_dataout[30]),
      .A2F_R_7_2(m0_m0_dataout[29]),
      .A2F_R_7_3(m0_m0_dataout[28]),
      .A2F_R_7_4(m0_m0_dataout[27]),
      .A2F_R_7_5(m0_m0_dataout[26]),
      .A2F_R_8_0(m0_m0_dataout[25]),
      .A2F_R_8_1(m0_m0_dataout[24]),
      .A2F_R_8_2(m0_m0_dataout[23]),
      .A2F_R_8_3(m0_m0_dataout[22]),
      .A2F_R_8_4(m0_m0_dataout[21]),
      .A2F_R_8_5(m0_m0_dataout[20]),
      .A2F_R_8_6(m0_m0_dataout[19]),
      .A2F_R_8_7(m0_m0_dataout[18]),
      .A2F_R_9_0(m0_m0_dataout[17]),
      .A2F_R_9_1(m0_m0_dataout[16]),
      .A2F_R_9_2(m0_m0_dataout[15]),
      .A2F_R_9_3(m0_m0_dataout[14]),
      .A2F_R_9_4(m0_m0_dataout[13]),
      .A2F_R_9_5(m0_m0_dataout[12]),
      .A2Freg_B_11_0(1'b0),
      .A2Freg_B_13_0(1'b0),
      .A2Freg_B_15_0(1'b0),
      .A2Freg_B_17_0(1'b0),
      .A2Freg_B_19_0(1'b0),
      .A2Freg_B_1_0(1'b0),
      .A2Freg_B_21_0(1'b0),
      .A2Freg_B_23_0(1'b0),
      .A2Freg_B_25_0(1'b0),
      .A2Freg_B_27_0(1'b0),
      .A2Freg_B_29_0(1'b0),
      .A2Freg_B_31_0(1'b0),
      .A2Freg_B_3_0(1'b0),
      .A2Freg_B_5_0(1'b0),
      .A2Freg_B_7_0(1'b0),
      .A2Freg_B_9_0(1'b0),
      .A2Freg_L_11_0(1'b0),
      .A2Freg_L_13_0(1'b0),
      .A2Freg_L_15_0(1'b0),
      .A2Freg_L_17_0(1'b0),
      .A2Freg_L_19_0(1'b0),
      .A2Freg_L_1_0(1'b0),
      .A2Freg_L_21_0(1'b0),
      .A2Freg_L_23_0(1'b0),
      .A2Freg_L_25_0(1'b0),
      .A2Freg_L_27_0(1'b0),
      .A2Freg_L_29_0(1'b0),
      .A2Freg_L_31_0(1'b0),
      .A2Freg_L_3_0(1'b0),
      .A2Freg_L_5_0(1'b0),
      .A2Freg_L_7_0(1'b0),
      .A2Freg_L_9_0(1'b0),
      .A2Freg_T_11_0(1'b0),
      .A2Freg_T_13_0(1'b0),
      .A2Freg_T_15_0(1'b0),
      .A2Freg_T_17_0(1'b0),
      .A2Freg_T_19_0(1'b0),
      .A2Freg_T_1_0(1'b0),
      .A2Freg_T_21_0(1'b0),
      .A2Freg_T_23_0(1'b0),
      .A2Freg_T_25_0(1'b0),
      .A2Freg_T_27_0(1'b0),
      .A2Freg_T_29_0(1'b0),
      .A2Freg_T_31_0(1'b0),
      .A2Freg_T_3_0(1'b0),
      .A2Freg_T_5_0(1'b0),
      .A2Freg_T_7_0(1'b0),
      .A2Freg_T_9_0(1'b0),
      .A2Freg_R_11_0(1'b0),
      .A2Freg_R_13_0(1'b0),
      .A2Freg_R_15_0(1'b0),
      .A2Freg_R_17_0(1'b0),
      .A2Freg_R_19_0(1'b0),
      .A2Freg_R_1_0(1'b0),
      .A2Freg_R_21_0(1'b0),
      .A2Freg_R_23_0(1'b0),
      .A2Freg_R_25_0(1'b0),
      .A2Freg_R_27_0(1'b0),
      .A2Freg_R_29_0(1'b0),
      .A2Freg_R_31_0(1'b0),
      .A2Freg_R_3_0(1'b0),
      .A2Freg_R_5_0(1'b0),
      .A2Freg_R_7_0(1'b0),
      .A2Freg_R_9_0(1'b0),
      .BL_CLK(fcb_blclk),
      .BL_DIN_0_(fcb_bl_din[0]),
      .BL_DIN_10_(fcb_bl_din[10]),
      .BL_DIN_11_(fcb_bl_din[11]),
      .BL_DIN_12_(fcb_bl_din[12]),
      .BL_DIN_13_(fcb_bl_din[13]),
      .BL_DIN_14_(fcb_bl_din[14]),
      .BL_DIN_15_(fcb_bl_din[15]),
      .BL_DIN_16_(fcb_bl_din[16]),
      .BL_DIN_17_(fcb_bl_din[17]),
      .BL_DIN_18_(fcb_bl_din[18]),
      .BL_DIN_19_(fcb_bl_din[19]),
      .BL_DIN_1_(fcb_bl_din[1]),
      .BL_DIN_20_(fcb_bl_din[20]),
      .BL_DIN_21_(fcb_bl_din[21]),
      .BL_DIN_22_(fcb_bl_din[22]),
      .BL_DIN_23_(fcb_bl_din[23]),
      .BL_DIN_24_(fcb_bl_din[24]),
      .BL_DIN_25_(fcb_bl_din[25]),
      .BL_DIN_26_(fcb_bl_din[26]),
      .BL_DIN_27_(fcb_bl_din[27]),
      .BL_DIN_28_(fcb_bl_din[28]),
      .BL_DIN_29_(fcb_bl_din[29]),
      .BL_DIN_2_(fcb_bl_din[2]),
      .BL_DIN_30_(fcb_bl_din[30]),
      .BL_DIN_31_(fcb_bl_din[31]),
      .BL_DIN_3_(fcb_bl_din[3]),
      .BL_DIN_4_(fcb_bl_din[4]),
      .BL_DIN_5_(fcb_bl_din[5]),
      .BL_DIN_6_(fcb_bl_din[6]),
      .BL_DIN_7_(fcb_bl_din[7]),
      .BL_DIN_8_(fcb_bl_din[8]),
      .BL_DIN_9_(fcb_bl_din[9]),
      .BL_PWRGATE_0_(fcb_bl_pwrgate[0]),
      .BL_PWRGATE_1_(fcb_bl_pwrgate[1]),
      .BL_PWRGATE_2_(fcb_bl_pwrgate[2]),
      .BL_PWRGATE_3_(fcb_bl_pwrgate[3]),
      .CLOAD_DIN_SEL(fcb_cload_din_sel),
      .DIN_INT_L_ONLY(fcb_din_int_l_only),
      .DIN_INT_R_ONLY(fcb_din_int_r_only),
      .DIN_SLC_TB_INT(fcb_din_slc_tb_int),
      .FB_CFG_DONE(fcb_fb_cfg_done),
      .FB_ISO_ENB(fcb_fb_iso_enb),
      .FB_SPE_IN_0_(FB_SPE_IN[0]),
      .FB_SPE_IN_1_(FB_SPE_IN[1]),
      .FB_SPE_IN_2_(FB_SPE_IN[2]),
      .FB_SPE_IN_3_(FB_SPE_IN[3]),
      .ISO_EN_0_(fcb_iso_en[0]),
      .ISO_EN_1_(fcb_iso_en[1]),
      .ISO_EN_2_(fcb_iso_en[2]),
      .ISO_EN_3_(fcb_iso_en[3]),
      .MLATCH(MLATCH),
      .M_0_(M[0]),
      .M_1_(M[1]),
      .M_2_(M[2]),
      .M_3_(M[3]),
      .M_4_(M[4]),
      .M_5_(M[5]),
      .NB(NB),
      .PB(PB),
      .PCHG_B(fcb_pchg_b),
      .PI_PWR_0_(fcb_pi_pwr[0]),
      .PI_PWR_1_(fcb_pi_pwr[1]),
      .PI_PWR_2_(fcb_pi_pwr[2]),
      .PI_PWR_3_(fcb_pi_pwr[3]),
      .POR(POR),
      .PROG_0_(fcb_prog[0]),
      .PROG_1_(fcb_prog[1]),
      .PROG_2_(fcb_prog[2]),
      .PROG_3_(fcb_prog[3]),
      .PROG_IFX(fcb_prog_ifx),
      .PWR_GATE(fcb_pwr_gate),
      .RE(fcb_re),
      .STM(STM),
      .VLP_CLKDIS_0_(fcb_vlp_clkdis[0]),
      .VLP_CLKDIS_1_(fcb_vlp_clkdis[1]),
      .VLP_CLKDIS_2_(fcb_vlp_clkdis[2]),
      .VLP_CLKDIS_3_(fcb_vlp_clkdis[3]),
      .VLP_CLKDIS_IFX(fcb_vlp_clkdis_ifx),
      .VLP_PWRDIS_0_(fcb_vlp_pwrdis[0]),
      .VLP_PWRDIS_1_(fcb_vlp_pwrdis[1]),
      .VLP_PWRDIS_2_(fcb_vlp_pwrdis[2]),
      .VLP_PWRDIS_3_(fcb_vlp_pwrdis[3]),
      .VLP_PWRDIS_IFX(fcb_vlp_pwrdis_ifx),
      .VLP_SRDIS_0_(fcb_vlp_srdis[0]),
      .VLP_SRDIS_1_(fcb_vlp_srdis[1]),
      .VLP_SRDIS_2_(fcb_vlp_srdis[2]),
      .VLP_SRDIS_3_(fcb_vlp_srdis[3]),
      .VLP_SRDIS_IFX(fcb_vlp_srdis_ifx),
      .WE(fcb_we),
      .WE_INT(fcb_we_int),
      .WL_CLK(fcb_wlclk),
      .WL_CLOAD_SEL_0_(fcb_wl_cload_sel[0]),
      .WL_CLOAD_SEL_1_(fcb_wl_cload_sel[1]),
      .WL_CLOAD_SEL_2_(fcb_wl_cload_sel[2]),
      .WL_DIN_0_(fcb_wl_din[0]),
      .WL_DIN_1_(fcb_wl_din[1]),
      .WL_DIN_2_(fcb_wl_din[2]),
      .WL_DIN_3_(fcb_wl_din[3]),
      .WL_DIN_4_(fcb_wl_din[4]),
      .WL_DIN_5_(fcb_wl_din[5]),
      .WL_EN(fcb_wl_en),
      .WL_INT_DIN_SEL(fcb_wl_int_din_sel),
      .WL_PWRGATE_0_(fcb_wl_pwrgate[0]),
      .WL_PWRGATE_1_(fcb_wl_pwrgate[1]),
      .WL_RESETB(fcb_wl_resetb),
      .WL_SEL_0_(fcb_wl_sel[0]),
      .WL_SEL_1_(fcb_wl_sel[1]),
      .WL_SEL_2_(fcb_wl_sel[2]),
      .WL_SEL_3_(fcb_wl_sel[3]),
      .WL_SEL_TB_INT(fcb_wl_sel_tb_int),
      .F2A_B_10_0(m1_m0_coef_in[20]),
      .F2A_B_10_1(m1_m0_coef_in[19]),
      .F2A_B_10_10(m1_m0_coef_in[10]),
      .F2A_B_10_11(m1_m0_coef_in[9]),
      .F2A_B_10_12(m1_m0_coef_in[8]),
      .F2A_B_10_13(m1_m0_coef_in[7]),
      .F2A_B_10_14(m1_m0_coef_in[6]),
      .F2A_B_10_15(m1_m0_coef_in[5]),
      .F2A_B_10_16(m1_m0_coef_in[4]),
      .F2A_B_10_17(m1_m0_coef_in[3]),
      .F2A_B_10_2(m1_m0_coef_in[18]),
      .F2A_B_10_3(m1_m0_coef_in[17]),
      .F2A_B_10_4(m1_m0_coef_in[16]),
      .F2A_B_10_5(m1_m0_coef_in[15]),
      .F2A_B_10_6(m1_m0_coef_in[14]),
      .F2A_B_10_7(m1_m0_coef_in[13]),
      .F2A_B_10_8(m1_m0_coef_in[12]),
      .F2A_B_10_9(m1_m0_coef_in[11]),
      .F2A_B_11_0(m1_m0_coef_in[2]),
      .F2A_B_11_1(m1_m0_coef_in[1]),
      .F2A_B_11_10(m1_coef_wdata[28]),
      .F2A_B_11_11(m1_coef_wdata[27]),
      .F2A_B_11_2(m1_m0_coef_in[0]),
      .F2A_B_11_3(m1_m0_mode[1]),
      .F2A_B_11_4(m1_m0_mode[0]),
      .F2A_B_11_5(m1_m0_tc),
      .F2A_B_11_6(m1_m0_reset),
      .F2A_B_11_7(m1_coef_wdata[31]),
      .F2A_B_11_8(m1_coef_wdata[30]),
      .F2A_B_11_9(m1_coef_wdata[29]),
      .F2A_B_12_0(m1_coef_wdata[26]),
      .F2A_B_12_1(m1_coef_wdata[25]),
      .F2A_B_12_10(m1_coef_wdata[16]),
      .F2A_B_12_11(m1_coef_wdata[15]),
      .F2A_B_12_12(m1_coef_wdata[14]),
      .F2A_B_12_13(m1_coef_wdata[13]),
      .F2A_B_12_14(m1_coef_wdata[12]),
      .F2A_B_12_15(m1_coef_wdata[11]),
      .F2A_B_12_16(m1_coef_wdata[10]),
      .F2A_B_12_17(m1_coef_wdata[9]),
      .F2A_B_12_2(m1_coef_wdata[24]),
      .F2A_B_12_3(m1_coef_wdata[23]),
      .F2A_B_12_4(m1_coef_wdata[22]),
      .F2A_B_12_5(m1_coef_wdata[21]),
      .F2A_B_12_6(m1_coef_wdata[20]),
      .F2A_B_12_7(m1_coef_wdata[19]),
      .F2A_B_12_8(m1_coef_wdata[18]),
      .F2A_B_12_9(m1_coef_wdata[17]),
      .F2A_B_13_0(m1_coef_wclk_int),
      .F2A_B_13_1(m1_coef_wdata[8]),
      .F2A_B_13_10(m1_coef_waddr[11]),
      .F2A_B_13_11(m1_coef_waddr[10]),
      .F2A_B_13_2(m1_coef_wdata[7]),
      .F2A_B_13_3(m1_coef_wdata[6]),
      .F2A_B_13_4(m1_coef_wdata[5]),
      .F2A_B_13_5(m1_coef_wdata[4]),
      .F2A_B_13_6(m1_coef_wdata[3]),
      .F2A_B_13_7(m1_coef_wdata[2]),
      .F2A_B_13_8(m1_coef_wdata[1]),
      .F2A_B_13_9(m1_coef_wdata[0]),
      .F2A_B_14_0(m1_coef_waddr[9]),
      .F2A_B_14_1(m1_coef_waddr[8]),
      .F2A_B_14_10(m1_coef_we),
      .F2A_B_14_11(m1_coef_wdsel),
      .F2A_B_14_12(m1_coef_rmode[1]),
      .F2A_B_14_13(m1_coef_rmode[0]),
      .F2A_B_14_14(m1_coef_raddr[11]),
      .F2A_B_14_15(m1_coef_raddr[10]),
      .F2A_B_14_16(m1_coef_raddr[9]),
      .F2A_B_14_17(m1_coef_raddr[8]),
      .F2A_B_14_2(m1_coef_waddr[7]),
      .F2A_B_14_3(m1_coef_waddr[6]),
      .F2A_B_14_4(m1_coef_waddr[5]),
      .F2A_B_14_5(m1_coef_waddr[4]),
      .F2A_B_14_6(m1_coef_waddr[3]),
      .F2A_B_14_7(m1_coef_waddr[2]),
      .F2A_B_14_8(m1_coef_waddr[1]),
      .F2A_B_14_9(m1_coef_waddr[0]),
      .F2A_B_15_0(m1_coef_rclk_int),
      .F2A_B_15_1(m1_coef_raddr[7]),
      .F2A_B_15_10(m1_coef_wmode[0]),
      .F2A_B_15_11(),
      .F2A_B_15_2(m1_coef_raddr[6]),
      .F2A_B_15_3(m1_coef_raddr[5]),
      .F2A_B_15_4(m1_coef_raddr[4]),
      .F2A_B_15_5(m1_coef_raddr[3]),
      .F2A_B_15_6(m1_coef_raddr[2]),
      .F2A_B_15_7(m1_coef_raddr[1]),
      .F2A_B_15_8(m1_coef_raddr[0]),
      .F2A_B_15_9(m1_coef_wmode[1]),
      .F2A_B_16_0(),
      .F2A_B_16_1(),
      .F2A_B_16_10(),
      .F2A_B_16_11(),
      .F2A_B_16_12(),
      .F2A_B_16_13(),
      .F2A_B_16_17(),
      .F2A_B_16_2(),
      .F2A_B_16_3(),
      .F2A_B_16_4(),
      .F2A_B_16_5(),
      .F2A_B_16_6(),
      .F2A_B_16_7(),
      .F2A_B_16_8(),
      .F2A_B_16_9(),
      .F2A_B_17_0(),
      .F2A_B_17_1(),
      .F2A_B_17_10(),
      .F2A_B_17_11(),
      .F2A_B_17_2(),
      .F2A_B_17_3(),
      .F2A_B_17_4(),
      .F2A_B_17_5(),
      .F2A_B_17_6(),
      .F2A_B_17_7(),
      .F2A_B_17_8(),
      .F2A_B_17_9(),
      .F2A_B_18_0(),
      .F2A_B_18_1(),
      .F2A_B_18_10(m1_m1_outsel[2]),
      .F2A_B_18_11(m1_m1_outsel[1]),
      .F2A_B_18_12(m1_m1_outsel[0]),
      .F2A_B_18_13(m1_m1_sat),
      .F2A_B_18_14(m1_m1_rnd),
      .F2A_B_18_15(m1_m1_clr),
      .F2A_B_18_16(m1_m1_clken),
      .F2A_B_18_17(),
      .F2A_B_18_2(),
      .F2A_B_18_3(),
      .F2A_B_18_4(),
      .F2A_B_18_5(),
      .F2A_B_18_6(),
      .F2A_B_18_7(m1_m1_outsel[5]),
      .F2A_B_18_8(m1_m1_outsel[4]),
      .F2A_B_18_9(m1_m1_outsel[3]),
      .F2A_B_19_0(m1_m1_clk_int),
      .F2A_B_19_1(m1_m1_osel),
      .F2A_B_19_10(m1_m1_coef_in[25]),
      .F2A_B_19_11(m1_m1_coef_in[24]),
      .F2A_B_19_2(m1_m1_tc),
      .F2A_B_19_3(m1_m1_reset),
      .F2A_B_19_4(m1_m1_coef_in[31]),
      .F2A_B_19_5(m1_m1_coef_in[30]),
      .F2A_B_19_6(m1_m1_coef_in[29]),
      .F2A_B_19_7(m1_m1_coef_in[28]),
      .F2A_B_19_8(m1_m1_coef_in[27]),
      .F2A_B_19_9(m1_m1_coef_in[26]),
      .F2A_B_1_0(),
      .F2A_B_1_1(),
      .F2A_B_1_10(),
      .F2A_B_1_11(),
      .F2A_B_1_2(),
      .F2A_B_1_3(),
      .F2A_B_1_4(),
      .F2A_B_1_5(),
      .F2A_B_1_6(),
      .F2A_B_1_7(),
      .F2A_B_1_8(),
      .F2A_B_1_9(),
      .F2A_B_20_0(m1_m1_coef_in[23]),
      .F2A_B_20_1(m1_m1_coef_in[22]),
      .F2A_B_20_10(m1_m1_coef_in[13]),
      .F2A_B_20_11(m1_m1_coef_in[12]),
      .F2A_B_20_12(m1_m1_coef_in[11]),
      .F2A_B_20_13(m1_m1_coef_in[10]),
      .F2A_B_20_14(m1_m1_coef_in[9]),
      .F2A_B_20_15(m1_m1_coef_in[8]),
      .F2A_B_20_16(m1_m1_coef_in[7]),
      .F2A_B_20_17(m1_m1_coef_in[6]),
      .F2A_B_20_2(m1_m1_coef_in[21]),
      .F2A_B_20_3(m1_m1_coef_in[20]),
      .F2A_B_20_4(m1_m1_coef_in[19]),
      .F2A_B_20_5(m1_m1_coef_in[18]),
      .F2A_B_20_6(m1_m1_coef_in[17]),
      .F2A_B_20_7(m1_m1_coef_in[16]),
      .F2A_B_20_8(m1_m1_coef_in[15]),
      .F2A_B_20_9(m1_m1_coef_in[14]),
      .F2A_B_21_0(m1_m1_coef_in[5]),
      .F2A_B_21_1(m1_m1_coef_in[4]),
      .F2A_B_21_10(m1_m1_oper_in[30]),
      .F2A_B_21_11(m1_m1_oper_in[29]),
      .F2A_B_21_2(m1_m1_coef_in[3]),
      .F2A_B_21_3(m1_m1_coef_in[2]),
      .F2A_B_21_4(m1_m1_coef_in[1]),
      .F2A_B_21_5(m1_m1_coef_in[0]),
      .F2A_B_21_6(m1_m1_mode[1]),
      .F2A_B_21_7(m1_m1_csel),
      .F2A_B_21_8(m1_m1_mode[0]),
      .F2A_B_21_9(m1_m1_oper_in[31]),
      .F2A_B_22_0(m1_m1_oper_in[28]),
      .F2A_B_22_1(m1_m1_oper_in[27]),
      .F2A_B_22_10(m1_m1_oper_in[18]),
      .F2A_B_22_11(m1_m1_oper_in[17]),
      .F2A_B_22_12(m1_m1_oper_in[16]),
      .F2A_B_22_13(m1_m1_oper_in[15]),
      .F2A_B_22_14(m1_m1_oper_in[14]),
      .F2A_B_22_15(m1_m1_oper_in[13]),
      .F2A_B_22_16(m1_m1_oper_in[12]),
      .F2A_B_22_17(m1_m1_oper_in[11]),
      .F2A_B_22_2(m1_m1_oper_in[26]),
      .F2A_B_22_3(m1_m1_oper_in[25]),
      .F2A_B_22_4(m1_m1_oper_in[24]),
      .F2A_B_22_5(m1_m1_oper_in[23]),
      .F2A_B_22_6(m1_m1_oper_in[22]),
      .F2A_B_22_7(m1_m1_oper_in[21]),
      .F2A_B_22_8(m1_m1_oper_in[20]),
      .F2A_B_22_9(m1_m1_oper_in[19]),
      .F2A_B_23_0(m1_m1_oper_in[10]),
      .F2A_B_23_1(m1_m1_oper_in[9]),
      .F2A_B_23_10(m1_m1_oper_in[0]),
      .F2A_B_23_11(),
      .F2A_B_23_2(m1_m1_oper_in[8]),
      .F2A_B_23_3(m1_m1_oper_in[7]),
      .F2A_B_23_4(m1_m1_oper_in[6]),
      .F2A_B_23_5(m1_m1_oper_in[5]),
      .F2A_B_23_6(m1_m1_oper_in[4]),
      .F2A_B_23_7(m1_m1_oper_in[3]),
      .F2A_B_23_8(m1_m1_oper_in[2]),
      .F2A_B_23_9(m1_m1_oper_in[1]),
      .F2A_B_24_0(),
      .F2A_B_24_1(),
      .F2A_B_24_10(),
      .F2A_B_24_11(),
      .F2A_B_24_12(),
      .F2A_B_24_13(),
      .F2A_B_24_14(),
      .F2A_B_24_15(),
      .F2A_B_24_16(m1_oper1_wdata[31]),
      .F2A_B_24_17(m1_oper1_wdata[30]),
      .F2A_B_24_2(),
      .F2A_B_24_3(),
      .F2A_B_24_4(),
      .F2A_B_24_5(),
      .F2A_B_24_6(),
      .F2A_B_24_7(),
      .F2A_B_24_8(),
      .F2A_B_24_9(),
      .F2A_B_25_0(m1_oper1_wdata[29]),
      .F2A_B_25_1(m1_oper1_wdata[28]),
      .F2A_B_25_10(m1_oper1_wdata[19]),
      .F2A_B_25_11(m1_oper1_wdata[18]),
      .F2A_B_25_2(m1_oper1_wdata[27]),
      .F2A_B_25_3(m1_oper1_wdata[26]),
      .F2A_B_25_4(m1_oper1_wdata[25]),
      .F2A_B_25_5(m1_oper1_wdata[24]),
      .F2A_B_25_6(m1_oper1_wdata[23]),
      .F2A_B_25_7(m1_oper1_wdata[22]),
      .F2A_B_25_8(m1_oper1_wdata[21]),
      .F2A_B_25_9(m1_oper1_wdata[20]),
      .F2A_B_26_0(m1_oper1_wdata[17]),
      .F2A_B_26_1(m1_oper1_wdata[16]),
      .F2A_B_26_10(m1_oper1_wdata[7]),
      .F2A_B_26_11(m1_oper1_wdata[6]),
      .F2A_B_26_12(m1_oper1_wdata[5]),
      .F2A_B_26_13(m1_oper1_wdata[4]),
      .F2A_B_26_14(m1_oper1_wdata[3]),
      .F2A_B_26_15(m1_oper1_wdata[2]),
      .F2A_B_26_16(m1_oper1_wdata[1]),
      .F2A_B_26_17(m1_oper1_wdata[0]),
      .F2A_B_26_2(m1_oper1_wdata[15]),
      .F2A_B_26_3(m1_oper1_wdata[14]),
      .F2A_B_26_4(m1_oper1_wdata[13]),
      .F2A_B_26_5(m1_oper1_wdata[12]),
      .F2A_B_26_6(m1_oper1_wdata[11]),
      .F2A_B_26_7(m1_oper1_wdata[10]),
      .F2A_B_26_8(m1_oper1_wdata[9]),
      .F2A_B_26_9(m1_oper1_wdata[8]),
      .F2A_B_27_0(m1_oper1_waddr[11]),
      .F2A_B_27_1(m1_oper1_waddr[10]),
      .F2A_B_27_10(m1_oper1_waddr[1]),
      .F2A_B_27_11(m1_oper1_waddr[0]),
      .F2A_B_27_2(m1_oper1_waddr[9]),
      .F2A_B_27_3(m1_oper1_waddr[8]),
      .F2A_B_27_4(m1_oper1_waddr[7]),
      .F2A_B_27_5(m1_oper1_waddr[6]),
      .F2A_B_27_6(m1_oper1_waddr[5]),
      .F2A_B_27_7(m1_oper1_waddr[4]),
      .F2A_B_27_8(m1_oper1_waddr[3]),
      .F2A_B_27_9(m1_oper1_waddr[2]),
      .F2A_B_28_0(m1_oper1_wclk_int),
      .F2A_B_28_1(m1_oper1_wmode[1]),
      .F2A_B_28_10(),
      .F2A_B_28_11(),
      .F2A_B_28_12(),
      .F2A_B_28_13(),
      .F2A_B_28_14(),
      .F2A_B_28_15(m1_oper1_rmode[1]),
      .F2A_B_28_16(m1_oper1_rmode[0]),
      .F2A_B_28_17(m1_oper1_raddr[11]),
      .F2A_B_28_2(m1_oper1_wmode[0]),
      .F2A_B_28_3(m1_oper1_wdsel),
      .F2A_B_28_4(m1_oper1_we),
      .F2A_B_28_5(),
      .F2A_B_28_6(),
      .F2A_B_28_7(),
      .F2A_B_28_8(),
      .F2A_B_28_9(),
      .F2A_B_29_0(m1_oper1_rclk_int),
      .F2A_B_29_1(m1_oper1_raddr[10]),
      .F2A_B_29_10(m1_oper1_raddr[1]),
      .F2A_B_29_11(m1_oper1_raddr[0]),
      .F2A_B_29_2(m1_oper1_raddr[9]),
      .F2A_B_29_3(m1_oper1_raddr[8]),
      .F2A_B_29_4(m1_oper1_raddr[7]),
      .F2A_B_29_5(m1_oper1_raddr[6]),
      .F2A_B_29_6(m1_oper1_raddr[5]),
      .F2A_B_29_7(m1_oper1_raddr[4]),
      .F2A_B_29_8(m1_oper1_raddr[3]),
      .F2A_B_29_9(m1_oper1_raddr[2]),
      .F2A_B_2_0(m1_oper0_wclk_int),
      .F2A_B_2_1(m1_oper0_wmode[1]),
      .F2A_B_2_10(m1_oper0_wdata[27]),
      .F2A_B_2_11(m1_oper0_wdata[26]),
      .F2A_B_2_12(m1_oper0_wdata[25]),
      .F2A_B_2_13(m1_oper0_wdata[24]),
      .F2A_B_2_14(m1_oper0_wdata[23]),
      .F2A_B_2_15(m1_oper0_wdata[22]),
      .F2A_B_2_16(m1_oper0_wdata[21]),
      .F2A_B_2_17(m1_oper0_wdata[20]),
      .F2A_B_2_2(m1_oper0_wmode[0]),
      .F2A_B_2_3(m1_oper0_wdsel),
      .F2A_B_2_4(m1_oper0_rmode[1]),
      .F2A_B_2_5(m1_oper0_rmode[0]),
      .F2A_B_2_6(m1_oper0_wdata[31]),
      .F2A_B_2_7(m1_oper0_wdata[30]),
      .F2A_B_2_8(m1_oper0_wdata[29]),
      .F2A_B_2_9(m1_oper0_wdata[28]),
      .F2A_B_30_0(),
      .F2A_B_30_1(),
      .F2A_B_30_10(),
      .F2A_B_30_11(),
      .F2A_B_30_12(),
      .F2A_B_30_13(),
      .F2A_B_30_14(),
      .F2A_B_30_15(),
      .F2A_B_30_16(),
      .F2A_B_30_17(),
      .F2A_B_30_2(),
      .F2A_B_30_3(),
      .F2A_B_30_4(),
      .F2A_B_30_5(),
      .F2A_B_30_6(),
      .F2A_B_30_7(),
      .F2A_B_30_8(),
      .F2A_B_30_9(),
      .F2A_B_31_0(),
      .F2A_B_31_1(),
      .F2A_B_31_10(),
      .F2A_B_31_11(),
      .F2A_B_31_2(),
      .F2A_B_31_3(),
      .F2A_B_31_4(),
      .F2A_B_31_5(),
      .F2A_B_31_6(),
      .F2A_B_31_7(),
      .F2A_B_31_8(),
      .F2A_B_31_9(),
      .F2A_B_32_0(),
      .F2A_B_32_1(),
      .F2A_B_32_10(),
      .F2A_B_32_11(),
      .F2A_B_32_12(),
      .F2A_B_32_13(),
      .F2A_B_32_14(),
      .F2A_B_32_15(),
      .F2A_B_32_16(),
      .F2A_B_32_17(),
      .F2A_B_32_2(),
      .F2A_B_32_3(),
      .F2A_B_32_4(),
      .F2A_B_32_5(),
      .F2A_B_32_6(),
      .F2A_B_32_7(),
      .F2A_B_32_8(),
      .F2A_B_32_9(),
      .F2A_B_3_0(m1_oper0_wdata[19]),
      .F2A_B_3_1(m1_oper0_wdata[18]),
      .F2A_B_3_10(m1_oper0_wdata[9]),
      .F2A_B_3_11(m1_oper0_wdata[8]),
      .F2A_B_3_2(m1_oper0_wdata[17]),
      .F2A_B_3_3(m1_oper0_wdata[16]),
      .F2A_B_3_4(m1_oper0_wdata[15]),
      .F2A_B_3_5(m1_oper0_wdata[14]),
      .F2A_B_3_6(m1_oper0_wdata[13]),
      .F2A_B_3_7(m1_oper0_wdata[12]),
      .F2A_B_3_8(m1_oper0_wdata[11]),
      .F2A_B_3_9(m1_oper0_wdata[10]),
      .F2A_B_4_0(m1_oper0_wdata[7]),
      .F2A_B_4_1(m1_oper0_wdata[6]),
      .F2A_B_4_10(m1_oper0_waddr[9]),
      .F2A_B_4_11(m1_oper0_waddr[8]),
      .F2A_B_4_12(m1_oper0_waddr[7]),
      .F2A_B_4_13(m1_oper0_waddr[6]),
      .F2A_B_4_14(m1_oper0_waddr[5]),
      .F2A_B_4_15(m1_oper0_waddr[4]),
      .F2A_B_4_16(m1_oper0_waddr[3]),
      .F2A_B_4_17(m1_oper0_waddr[2]),
      .F2A_B_4_2(m1_oper0_wdata[5]),
      .F2A_B_4_3(m1_oper0_wdata[4]),
      .F2A_B_4_4(m1_oper0_wdata[3]),
      .F2A_B_4_5(m1_oper0_wdata[2]),
      .F2A_B_4_6(m1_oper0_wdata[1]),
      .F2A_B_4_7(m1_oper0_wdata[0]),
      .F2A_B_4_8(m1_oper0_waddr[11]),
      .F2A_B_4_9(m1_oper0_waddr[10]),
      .F2A_B_5_0(m1_oper0_waddr[1]),
      .F2A_B_5_1(m1_oper0_waddr[0]),
      .F2A_B_5_10(m1_oper0_raddr[4]),
      .F2A_B_5_11(m1_oper0_raddr[3]),
      .F2A_B_5_2(m1_oper0_we),
      .F2A_B_5_3(m1_oper0_raddr[11]),
      .F2A_B_5_4(m1_oper0_raddr[10]),
      .F2A_B_5_5(m1_oper0_raddr[9]),
      .F2A_B_5_6(m1_oper0_raddr[8]),
      .F2A_B_5_7(m1_oper0_raddr[7]),
      .F2A_B_5_8(m1_oper0_raddr[6]),
      .F2A_B_5_9(m1_oper0_raddr[5]),
      .F2A_B_6_0(m1_oper0_rclk_int),
      .F2A_B_6_1(m1_oper0_raddr[2]),
      .F2A_B_6_10(m1_m0_outsel[1]),
      .F2A_B_6_11(m1_m0_outsel[0]),
      .F2A_B_6_12(m1_m0_sat),
      .F2A_B_6_13(m1_m0_rnd),
      .F2A_B_6_14(m1_m0_clr),
      .F2A_B_6_15(m1_m0_oper_in[31]),
      .F2A_B_6_16(m1_m0_oper_in[30]),
      .F2A_B_6_17(m1_m0_oper_in[29]),
      .F2A_B_6_2(m1_oper0_raddr[1]),
      .F2A_B_6_3(m1_oper0_raddr[0]),
      .F2A_B_6_4(m1_m0_osel),
      .F2A_B_6_5(m1_m0_clken),
      .F2A_B_6_6(m1_m0_outsel[5]),
      .F2A_B_6_7(m1_m0_outsel[4]),
      .F2A_B_6_8(m1_m0_outsel[3]),
      .F2A_B_6_9(m1_m0_outsel[2]),
      .F2A_B_7_0(m1_m0_clk_int),
      .F2A_B_7_1(m1_m0_oper_in[28]),
      .F2A_B_7_10(m1_m0_oper_in[19]),
      .F2A_B_7_11(m1_m0_oper_in[18]),
      .F2A_B_7_2(m1_m0_oper_in[27]),
      .F2A_B_7_3(m1_m0_oper_in[26]),
      .F2A_B_7_4(m1_m0_oper_in[25]),
      .F2A_B_7_5(m1_m0_oper_in[24]),
      .F2A_B_7_6(m1_m0_oper_in[23]),
      .F2A_B_7_7(m1_m0_oper_in[22]),
      .F2A_B_7_8(m1_m0_oper_in[21]),
      .F2A_B_7_9(m1_m0_oper_in[20]),
      .F2A_B_8_0(m1_m0_oper_in[17]),
      .F2A_B_8_1(m1_m0_oper_in[16]),
      .F2A_B_8_10(m1_m0_oper_in[7]),
      .F2A_B_8_11(m1_m0_oper_in[6]),
      .F2A_B_8_12(m1_m0_oper_in[5]),
      .F2A_B_8_13(m1_m0_oper_in[4]),
      .F2A_B_8_14(m1_m0_oper_in[3]),
      .F2A_B_8_15(m1_m0_oper_in[2]),
      .F2A_B_8_16(m1_m0_oper_in[1]),
      .F2A_B_8_17(m1_m0_oper_in[0]),
      .F2A_B_8_2(m1_m0_oper_in[15]),
      .F2A_B_8_3(m1_m0_oper_in[14]),
      .F2A_B_8_4(m1_m0_oper_in[13]),
      .F2A_B_8_5(m1_m0_oper_in[12]),
      .F2A_B_8_6(m1_m0_oper_in[11]),
      .F2A_B_8_7(m1_m0_oper_in[10]),
      .F2A_B_8_8(m1_m0_oper_in[9]),
      .F2A_B_8_9(m1_m0_oper_in[8]),
      .F2A_B_9_0(m1_m0_csel),
      .F2A_B_9_1(m1_m0_coef_in[31]),
      .F2A_B_9_10(m1_m0_coef_in[22]),
      .F2A_B_9_11(m1_m0_coef_in[21]),
      .F2A_B_9_2(m1_m0_coef_in[30]),
      .F2A_B_9_3(m1_m0_coef_in[29]),
      .F2A_B_9_4(m1_m0_coef_in[28]),
      .F2A_B_9_5(m1_m0_coef_in[27]),
      .F2A_B_9_6(m1_m0_coef_in[26]),
      .F2A_B_9_7(m1_m0_coef_in[25]),
      .F2A_B_9_8(m1_m0_coef_in[24]),
      .F2A_B_9_9(m1_m0_coef_in[23]),
      .F2A_L_10_0(),
      .F2A_L_10_1(),
      .F2A_L_10_10(),
      .F2A_L_10_11(),
      .F2A_L_10_12(),
      .F2A_L_10_13(),
      .F2A_L_10_14(),
      .F2A_L_10_15(),
      .F2A_L_10_16(),
      .F2A_L_10_17(),
      .F2A_L_10_2(),
      .F2A_L_10_3(),
      .F2A_L_10_4(),
      .F2A_L_10_5(),
      .F2A_L_10_6(),
      .F2A_L_10_7(),
      .F2A_L_10_8(),
      .F2A_L_10_9(),
      .F2A_L_11_0(),
      .F2A_L_11_1(),
      .F2A_L_11_10(),
      .F2A_L_11_11(),
      .F2A_L_11_2(),
      .F2A_L_11_3(),
      .F2A_L_11_4(),
      .F2A_L_11_5(),
      .F2A_L_11_6(),
      .F2A_L_11_7(),
      .F2A_L_11_8(),
      .F2A_L_11_9(),
      .F2A_L_12_0(),
      .F2A_L_12_1(),
      .F2A_L_12_10(lint_RDATA[2]),
      .F2A_L_12_11(lint_RDATA[3]),
      .F2A_L_12_12(lint_RDATA[4]),
      .F2A_L_12_13(lint_RDATA[5]),
      .F2A_L_12_14(lint_RDATA[6]),
      .F2A_L_12_15(lint_RDATA[7]),
      .F2A_L_12_16(lint_RDATA[8]),
      .F2A_L_12_17(),
      .F2A_L_12_2(),
      .F2A_L_12_3(),
      .F2A_L_12_4(),
      .F2A_L_12_5(),
      .F2A_L_12_6(),
      .F2A_L_12_7(),
      .F2A_L_12_8(lint_RDATA[0]),
      .F2A_L_12_9(lint_RDATA[1]),
      .F2A_L_13_0(lint_RDATA[9]),
      .F2A_L_13_1(lint_RDATA[10]),
      .F2A_L_13_10(),
      .F2A_L_13_11(),
      .F2A_L_13_2(lint_RDATA[11]),
      .F2A_L_13_3(lint_RDATA[12]),
      .F2A_L_13_4(lint_RDATA[13]),
      .F2A_L_13_5(lint_RDATA[14]),
      .F2A_L_13_6(lint_RDATA[15]),
      .F2A_L_13_7(),
      .F2A_L_13_8(),
      .F2A_L_13_9(),
      .F2A_L_14_0(lint_clk_int),
      .F2A_L_14_1(lint_RDATA[16]),
      .F2A_L_14_10(),
      .F2A_L_14_11(),
      .F2A_L_14_12(),
      .F2A_L_14_13(),
      .F2A_L_14_14(),
      .F2A_L_14_15(),
      .F2A_L_14_16(),
      .F2A_L_14_17(),
      .F2A_L_14_2(lint_RDATA[17]),
      .F2A_L_14_3(lint_RDATA[18]),
      .F2A_L_14_4(lint_RDATA[19]),
      .F2A_L_14_5(lint_RDATA[20]),
      .F2A_L_14_6(lint_RDATA[21]),
      .F2A_L_14_7(lint_RDATA[22]),
      .F2A_L_14_8(lint_RDATA[23]),
      .F2A_L_14_9(lint_VALID),
      .F2A_L_15_0(lint_RDATA[24]),
      .F2A_L_15_1(lint_RDATA[25]),
      .F2A_L_15_10(),
      .F2A_L_15_11(),
      .F2A_L_15_2(lint_RDATA[26]),
      .F2A_L_15_3(lint_RDATA[27]),
      .F2A_L_15_4(lint_RDATA[28]),
      .F2A_L_15_5(lint_RDATA[29]),
      .F2A_L_15_6(lint_RDATA[30]),
      .F2A_L_15_7(lint_RDATA[31]),
      .F2A_L_15_8(lint_GNT),
      .F2A_L_15_9(),
      .F2A_L_16_0(),
      .F2A_L_16_1(),
      .F2A_L_16_10(),
      .F2A_L_16_11(),
      .F2A_L_16_12(),
      .F2A_L_16_13(),
      .F2A_L_16_14(),
      .F2A_L_16_15(),
      .F2A_L_16_16(),
      .F2A_L_16_17(),
      .F2A_L_16_2(),
      .F2A_L_16_3(),
      .F2A_L_16_4(),
      .F2A_L_16_5(),
      .F2A_L_16_6(),
      .F2A_L_16_7(),
      .F2A_L_16_8(),
      .F2A_L_16_9(),
      .F2A_L_17_0(fpgaio_out[64]),
      .F2A_L_17_1(fpgaio_oe[64]),
      .F2A_L_17_10(),
      .F2A_L_17_11(),
      .F2A_L_17_2(fpgaio_out[65]),
      .F2A_L_17_3(fpgaio_oe[65]),
      .F2A_L_17_4(fpgaio_out[66]),
      .F2A_L_17_5(fpgaio_oe[66]),
      .F2A_L_17_6(fpgaio_out[67]),
      .F2A_L_17_7(fpgaio_oe[67]),
      .F2A_L_17_8(),
      .F2A_L_17_9(),
      .F2A_L_18_0(fpgaio_out[68]),
      .F2A_L_18_1(fpgaio_oe[68]),
      .F2A_L_18_10(fpgaio_out[73]),
      .F2A_L_18_11(fpgaio_oe[73]),
      .F2A_L_18_12(fpgaio_out[74]),
      .F2A_L_18_13(fpgaio_oe[74]),
      .F2A_L_18_14(fpgaio_out[75]),
      .F2A_L_18_15(fpgaio_oe[75]),
      .F2A_L_18_16(),
      .F2A_L_18_17(),
      .F2A_L_18_2(fpgaio_out[69]),
      .F2A_L_18_3(fpgaio_oe[69]),
      .F2A_L_18_4(fpgaio_out[70]),
      .F2A_L_18_5(fpgaio_oe[70]),
      .F2A_L_18_6(fpgaio_out[71]),
      .F2A_L_18_7(fpgaio_oe[71]),
      .F2A_L_18_8(fpgaio_out[72]),
      .F2A_L_18_9(fpgaio_oe[72]),
      .F2A_L_19_0(fpgaio_out[76]),
      .F2A_L_19_1(fpgaio_oe[76]),
      .F2A_L_19_10(),
      .F2A_L_19_11(),
      .F2A_L_19_2(fpgaio_out[77]),
      .F2A_L_19_3(fpgaio_oe[77]),
      .F2A_L_19_4(fpgaio_out[78]),
      .F2A_L_19_5(fpgaio_oe[78]),
      .F2A_L_19_6(fpgaio_out[79]),
      .F2A_L_19_7(fpgaio_oe[79]),
      .F2A_L_19_8(),
      .F2A_L_19_9(),
      .F2A_L_1_0(),
      .F2A_L_1_1(),
      .F2A_L_1_10(),
      .F2A_L_1_11(),
      .F2A_L_1_2(),
      .F2A_L_1_3(),
      .F2A_L_1_4(),
      .F2A_L_1_5(),
      .F2A_L_1_6(),
      .F2A_L_1_7(),
      .F2A_L_1_8(),
      .F2A_L_1_9(),
      .F2A_L_20_0(status_out[0]),
      .F2A_L_20_1(status_out[1]),
      .F2A_L_20_10(status_out[10]),
      .F2A_L_20_11(status_out[11]),
      .F2A_L_20_12(status_out[12]),
      .F2A_L_20_13(status_out[13]),
      .F2A_L_20_14(status_out[14]),
      .F2A_L_20_15(status_out[15]),
      .F2A_L_20_16(status_out[16]),
      .F2A_L_20_17(status_out[17]),
      .F2A_L_20_2(status_out[2]),
      .F2A_L_20_3(status_out[3]),
      .F2A_L_20_4(status_out[4]),
      .F2A_L_20_5(status_out[5]),
      .F2A_L_20_6(status_out[6]),
      .F2A_L_20_7(status_out[7]),
      .F2A_L_20_8(status_out[8]),
      .F2A_L_20_9(status_out[9]),
      .F2A_L_21_0(status_out[18]),
      .F2A_L_21_1(status_out[19]),
      .F2A_L_21_10(status_out[28]),
      .F2A_L_21_11(status_out[29]),
      .F2A_L_21_2(status_out[20]),
      .F2A_L_21_3(status_out[21]),
      .F2A_L_21_4(status_out[22]),
      .F2A_L_21_5(status_out[23]),
      .F2A_L_21_6(status_out[24]),
      .F2A_L_21_7(status_out[25]),
      .F2A_L_21_8(status_out[26]),
      .F2A_L_21_9(status_out[27]),
      .F2A_L_22_0(status_out[30]),
      .F2A_L_22_1(status_out[31]),
      .F2A_L_22_10(),
      .F2A_L_22_11(),
      .F2A_L_22_12(),
      .F2A_L_22_13(),
      .F2A_L_22_14(),
      .F2A_L_22_15(),
      .F2A_L_22_16(),
      .F2A_L_22_17(),
      .F2A_L_22_2(),
      .F2A_L_22_3(),
      .F2A_L_22_4(),
      .F2A_L_22_5(),
      .F2A_L_22_6(),
      .F2A_L_22_7(),
      .F2A_L_22_8(),
      .F2A_L_22_9(),
      .F2A_L_23_0(),
      .F2A_L_23_1(),
      .F2A_L_23_10(),
      .F2A_L_23_11(),
      .F2A_L_23_2(),
      .F2A_L_23_3(),
      .F2A_L_23_4(),
      .F2A_L_23_5(),
      .F2A_L_23_6(),
      .F2A_L_23_7(),
      .F2A_L_23_8(),
      .F2A_L_23_9(),
      .F2A_L_24_0(),
      .F2A_L_24_1(),
      .F2A_L_24_10(),
      .F2A_L_24_11(),
      .F2A_L_24_12(),
      .F2A_L_24_13(),
      .F2A_L_24_14(),
      .F2A_L_24_15(),
      .F2A_L_24_16(),
      .F2A_L_24_17(),
      .F2A_L_24_2(),
      .F2A_L_24_3(),
      .F2A_L_24_4(),
      .F2A_L_24_5(),
      .F2A_L_24_6(),
      .F2A_L_24_7(),
      .F2A_L_24_8(),
      .F2A_L_24_9(),
      .F2A_L_25_0(fpgaio_out[32]),
      .F2A_L_25_1(fpgaio_oe[32]),
      .F2A_L_25_10(),
      .F2A_L_25_11(),
      .F2A_L_25_2(fpgaio_out[33]),
      .F2A_L_25_3(fpgaio_oe[33]),
      .F2A_L_25_4(fpgaio_out[34]),
      .F2A_L_25_5(fpgaio_oe[34]),
      .F2A_L_25_6(fpgaio_out[35]),
      .F2A_L_25_7(fpgaio_oe[35]),
      .F2A_L_25_8(events_o[8]),
      .F2A_L_25_9(),
      .F2A_L_26_0(fpgaio_out[36]),
      .F2A_L_26_1(fpgaio_oe[36]),
      .F2A_L_26_10(),
      .F2A_L_26_11(),
      .F2A_L_26_12(),
      .F2A_L_26_13(),
      .F2A_L_26_14(),
      .F2A_L_26_15(),
      .F2A_L_26_16(),
      .F2A_L_26_17(),
      .F2A_L_26_2(fpgaio_out[37]),
      .F2A_L_26_3(fpgaio_oe[37]),
      .F2A_L_26_4(fpgaio_out[38]),
      .F2A_L_26_5(fpgaio_oe[38]),
      .F2A_L_26_6(fpgaio_out[39]),
      .F2A_L_26_7(fpgaio_oe[39]),
      .F2A_L_26_8(events_o[9]),
      .F2A_L_26_9(),
      .F2A_L_27_0(fpgaio_out[40]),
      .F2A_L_27_1(fpgaio_oe[40]),
      .F2A_L_27_10(),
      .F2A_L_27_11(),
      .F2A_L_27_2(fpgaio_out[41]),
      .F2A_L_27_3(fpgaio_oe[41]),
      .F2A_L_27_4(fpgaio_out[42]),
      .F2A_L_27_5(fpgaio_oe[42]),
      .F2A_L_27_6(fpgaio_out[43]),
      .F2A_L_27_7(fpgaio_oe[43]),
      .F2A_L_27_8(events_o[10]),
      .F2A_L_27_9(),
      .F2A_L_28_0(fpgaio_out[44]),
      .F2A_L_28_1(fpgaio_oe[44]),
      .F2A_L_28_10(),
      .F2A_L_28_11(),
      .F2A_L_28_12(),
      .F2A_L_28_13(),
      .F2A_L_28_14(),
      .F2A_L_28_15(),
      .F2A_L_28_16(),
      .F2A_L_28_17(),
      .F2A_L_28_2(fpgaio_out[45]),
      .F2A_L_28_3(fpgaio_oe[45]),
      .F2A_L_28_4(fpgaio_out[46]),
      .F2A_L_28_5(fpgaio_oe[46]),
      .F2A_L_28_6(fpgaio_out[47]),
      .F2A_L_28_7(fpgaio_oe[47]),
      .F2A_L_28_8(events_o[11]),
      .F2A_L_28_9(),
      .F2A_L_29_0(fpgaio_out[48]),
      .F2A_L_29_1(fpgaio_oe[48]),
      .F2A_L_29_10(),
      .F2A_L_29_11(),
      .F2A_L_29_2(fpgaio_out[49]),
      .F2A_L_29_3(fpgaio_oe[49]),
      .F2A_L_29_4(fpgaio_out[50]),
      .F2A_L_29_5(fpgaio_oe[50]),
      .F2A_L_29_6(fpgaio_out[51]),
      .F2A_L_29_7(fpgaio_oe[51]),
      .F2A_L_29_8(events_o[12]),
      .F2A_L_29_9(),
      .F2A_L_2_0(fpgaio_out[0]),
      .F2A_L_2_1(fpgaio_oe[0]),
      .F2A_L_2_10(),
      .F2A_L_2_11(),
      .F2A_L_2_12(),
      .F2A_L_2_13(),
      .F2A_L_2_14(),
      .F2A_L_2_15(),
      .F2A_L_2_16(),
      .F2A_L_2_17(),
      .F2A_L_2_2(fpgaio_out[1]),
      .F2A_L_2_3(fpgaio_oe[1]),
      .F2A_L_2_4(fpgaio_out[2]),
      .F2A_L_2_5(fpgaio_oe[2]),
      .F2A_L_2_6(fpgaio_out[3]),
      .F2A_L_2_7(fpgaio_oe[3]),
      .F2A_L_2_8(events_o[0]),
      .F2A_L_2_9(),
      .F2A_L_30_0(fpgaio_out[52]),
      .F2A_L_30_1(fpgaio_oe[52]),
      .F2A_L_30_10(),
      .F2A_L_30_11(),
      .F2A_L_30_12(),
      .F2A_L_30_13(),
      .F2A_L_30_14(),
      .F2A_L_30_15(),
      .F2A_L_30_16(),
      .F2A_L_30_17(),
      .F2A_L_30_2(fpgaio_out[53]),
      .F2A_L_30_3(fpgaio_oe[53]),
      .F2A_L_30_4(fpgaio_out[54]),
      .F2A_L_30_5(fpgaio_oe[54]),
      .F2A_L_30_6(fpgaio_out[55]),
      .F2A_L_30_7(fpgaio_oe[55]),
      .F2A_L_30_8(events_o[13]),
      .F2A_L_30_9(),
      .F2A_L_31_0(fpgaio_out[56]),
      .F2A_L_31_1(fpgaio_oe[56]),
      .F2A_L_31_10(),
      .F2A_L_31_11(),
      .F2A_L_31_2(fpgaio_out[57]),
      .F2A_L_31_3(fpgaio_oe[57]),
      .F2A_L_31_4(fpgaio_out[58]),
      .F2A_L_31_5(fpgaio_oe[58]),
      .F2A_L_31_6(fpgaio_out[59]),
      .F2A_L_31_7(fpgaio_oe[59]),
      .F2A_L_31_8(events_o[14]),
      .F2A_L_31_9(),
      .F2A_L_32_0(fpgaio_out[60]),
      .F2A_L_32_1(fpgaio_oe[60]),
      .F2A_L_32_10(),
      .F2A_L_32_11(),
      .F2A_L_32_12(),
      .F2A_L_32_13(),
      .F2A_L_32_14(),
      .F2A_L_32_15(),
      .F2A_L_32_16(),
      .F2A_L_32_17(),
      .F2A_L_32_2(fpgaio_out[61]),
      .F2A_L_32_3(fpgaio_oe[61]),
      .F2A_L_32_4(fpgaio_out[62]),
      .F2A_L_32_5(fpgaio_oe[62]),
      .F2A_L_32_6(fpgaio_out[63]),
      .F2A_L_32_7(fpgaio_oe[63]),
      .F2A_L_32_8(events_o[15]),
      .F2A_L_32_9(),
      .F2A_L_3_0(fpgaio_out[4]),
      .F2A_L_3_1(fpgaio_oe[4]),
      .F2A_L_3_10(),
      .F2A_L_3_11(),
      .F2A_L_3_2(fpgaio_out[5]),
      .F2A_L_3_3(fpgaio_oe[5]),
      .F2A_L_3_4(fpgaio_out[6]),
      .F2A_L_3_5(fpgaio_oe[6]),
      .F2A_L_3_6(fpgaio_out[7]),
      .F2A_L_3_7(fpgaio_oe[7]),
      .F2A_L_3_8(events_o[1]),
      .F2A_L_3_9(),
      .F2A_L_4_0(fpgaio_out[8]),
      .F2A_L_4_1(fpgaio_oe[8]),
      .F2A_L_4_10(fpgaio_oe[12]),
      .F2A_L_4_11(fpgaio_out[13]),
      .F2A_L_4_12(fpgaio_oe[13]),
      .F2A_L_4_13(fpgaio_out[14]),
      .F2A_L_4_14(fpgaio_oe[14]),
      .F2A_L_4_15(),
      .F2A_L_4_16(),
      .F2A_L_4_17(),
      .F2A_L_4_2(fpgaio_out[9]),
      .F2A_L_4_3(fpgaio_oe[9]),
      .F2A_L_4_4(fpgaio_out[10]),
      .F2A_L_4_5(fpgaio_oe[10]),
      .F2A_L_4_6(fpgaio_out[11]),
      .F2A_L_4_7(fpgaio_oe[11]),
      .F2A_L_4_8(events_o[2]),
      .F2A_L_4_9(fpgaio_out[12]),
      .F2A_L_5_0(fpgaio_out[15]),
      .F2A_L_5_1(fpgaio_oe[15]),
      .F2A_L_5_10(fpgaio_oe[19]),
      .F2A_L_5_11(events_o[4]),
      .F2A_L_5_2(events_o[3]),
      .F2A_L_5_3(fpgaio_out[16]),
      .F2A_L_5_4(fpgaio_oe[16]),
      .F2A_L_5_5(fpgaio_out[17]),
      .F2A_L_5_6(fpgaio_oe[17]),
      .F2A_L_5_7(fpgaio_out[18]),
      .F2A_L_5_8(fpgaio_oe[18]),
      .F2A_L_5_9(fpgaio_out[19]),
      .F2A_L_6_0(fpgaio_out[20]),
      .F2A_L_6_1(fpgaio_oe[20]),
      .F2A_L_6_10(fpgaio_oe[24]),
      .F2A_L_6_11(fpgaio_out[25]),
      .F2A_L_6_12(fpgaio_oe[25]),
      .F2A_L_6_13(fpgaio_out[26]),
      .F2A_L_6_14(fpgaio_oe[26]),
      .F2A_L_6_15(fpgaio_out[27]),
      .F2A_L_6_16(fpgaio_oe[27]),
      .F2A_L_6_17(events_o[6]),
      .F2A_L_6_2(fpgaio_out[21]),
      .F2A_L_6_3(fpgaio_oe[21]),
      .F2A_L_6_4(fpgaio_out[22]),
      .F2A_L_6_5(fpgaio_oe[22]),
      .F2A_L_6_6(fpgaio_out[23]),
      .F2A_L_6_7(fpgaio_oe[23]),
      .F2A_L_6_8(events_o[5]),
      .F2A_L_6_9(fpgaio_out[24]),
      .F2A_L_7_0(),
      .F2A_L_7_1(),
      .F2A_L_7_10(),
      .F2A_L_7_11(),
      .F2A_L_7_2(),
      .F2A_L_7_3(),
      .F2A_L_7_4(),
      .F2A_L_7_5(),
      .F2A_L_7_6(),
      .F2A_L_7_7(),
      .F2A_L_7_8(),
      .F2A_L_7_9(),
      .F2A_L_8_0(fpgaio_out[28]),
      .F2A_L_8_1(fpgaio_oe[28]),
      .F2A_L_8_10(),
      .F2A_L_8_11(),
      .F2A_L_8_12(),
      .F2A_L_8_13(),
      .F2A_L_8_14(),
      .F2A_L_8_15(),
      .F2A_L_8_16(),
      .F2A_L_8_17(),
      .F2A_L_8_2(fpgaio_out[29]),
      .F2A_L_8_3(fpgaio_oe[29]),
      .F2A_L_8_4(fpgaio_out[30]),
      .F2A_L_8_5(fpgaio_oe[30]),
      .F2A_L_8_6(fpgaio_out[31]),
      .F2A_L_8_7(fpgaio_oe[31]),
      .F2A_L_8_8(events_o[7]),
      .F2A_L_8_9(),
      .F2A_L_9_0(),
      .F2A_L_9_1(),
      .F2A_L_9_10(),
      .F2A_L_9_11(),
      .F2A_L_9_2(),
      .F2A_L_9_3(),
      .F2A_L_9_4(),
      .F2A_L_9_5(),
      .F2A_L_9_6(),
      .F2A_L_9_7(),
      .F2A_L_9_8(),
      .F2A_L_9_9(),
      .F2A_T_10_0(tcdm_wdata_p1[0]),
      .F2A_T_10_1(tcdm_wdata_p1[1]),
      .F2A_T_10_10(tcdm_addr_p1[5]),
      .F2A_T_10_11(tcdm_addr_p1[6]),
      .F2A_T_10_12(tcdm_addr_p1[7]),
      .F2A_T_10_13(tcdm_addr_p1[8]),
      .F2A_T_10_14(tcdm_addr_p1[9]),
      .F2A_T_10_15(),
      .F2A_T_10_16(),
      .F2A_T_10_17(),
      .F2A_T_10_2(tcdm_wdata_p1[2]),
      .F2A_T_10_3(tcdm_wdata_p1[3]),
      .F2A_T_10_4(tcdm_wdata_p1[4]),
      .F2A_T_10_5(tcdm_wdata_p1[5]),
      .F2A_T_10_6(tcdm_wdata_p1[6]),
      .F2A_T_10_7(tcdm_wdata_p1[7]),
      .F2A_T_10_8(),
      .F2A_T_10_9(tcdm_addr_p1[4]),
      .F2A_T_11_0(tcdm_wdata_p1[8]),
      .F2A_T_11_1(tcdm_wdata_p1[9]),
      .F2A_T_11_10(tcdm_addr_p1[12]),
      .F2A_T_11_11(tcdm_addr_p1[13]),
      .F2A_T_11_2(tcdm_wdata_p1[10]),
      .F2A_T_11_3(tcdm_wdata_p1[11]),
      .F2A_T_11_4(tcdm_wdata_p1[12]),
      .F2A_T_11_5(tcdm_wdata_p1[13]),
      .F2A_T_11_6(tcdm_wdata_p1[14]),
      .F2A_T_11_7(tcdm_wdata_p1[15]),
      .F2A_T_11_8(tcdm_addr_p1[10]),
      .F2A_T_11_9(tcdm_addr_p1[11]),
      .F2A_T_12_0(tcdm_wdata_p1[16]),
      .F2A_T_12_1(tcdm_wdata_p1[17]),
      .F2A_T_12_10(),
      .F2A_T_12_11(),
      .F2A_T_12_12(tcdm_addr_p1[14]),
      .F2A_T_12_13(tcdm_addr_p1[15]),
      .F2A_T_12_14(tcdm_addr_p1[16]),
      .F2A_T_12_15(tcdm_addr_p1[17]),
      .F2A_T_12_16(tcdm_addr_p1[18]),
      .F2A_T_12_17(tcdm_addr_p1[19]),
      .F2A_T_12_2(tcdm_wdata_p1[18]),
      .F2A_T_12_3(tcdm_wdata_p1[19]),
      .F2A_T_12_4(tcdm_wdata_p1[20]),
      .F2A_T_12_5(tcdm_wdata_p1[21]),
      .F2A_T_12_6(tcdm_wdata_p1[22]),
      .F2A_T_12_7(tcdm_wdata_p1[23]),
      .F2A_T_12_8(),
      .F2A_T_12_9(),
      .F2A_T_13_0(tcdm_wdata_p1[24]),
      .F2A_T_13_1(tcdm_wdata_p1[25]),
      .F2A_T_13_10(),
      .F2A_T_13_11(),
      .F2A_T_13_2(tcdm_wdata_p1[26]),
      .F2A_T_13_3(tcdm_wdata_p1[27]),
      .F2A_T_13_4(tcdm_wdata_p1[28]),
      .F2A_T_13_5(tcdm_wdata_p1[29]),
      .F2A_T_13_6(tcdm_wdata_p1[30]),
      .F2A_T_13_7(tcdm_wdata_p1[31]),
      .F2A_T_13_8(),
      .F2A_T_13_9(),
      .F2A_T_14_0(),
      .F2A_T_14_1(),
      .F2A_T_14_10(),
      .F2A_T_14_11(),
      .F2A_T_14_12(),
      .F2A_T_14_13(),
      .F2A_T_14_14(),
      .F2A_T_14_15(),
      .F2A_T_14_16(),
      .F2A_T_14_17(),
      .F2A_T_14_2(),
      .F2A_T_14_3(),
      .F2A_T_14_4(),
      .F2A_T_14_5(),
      .F2A_T_14_6(),
      .F2A_T_14_7(),
      .F2A_T_14_8(),
      .F2A_T_14_9(),
      .F2A_T_15_0(),
      .F2A_T_15_1(),
      .F2A_T_15_10(),
      .F2A_T_15_11(),
      .F2A_T_15_2(),
      .F2A_T_15_3(),
      .F2A_T_15_4(),
      .F2A_T_15_5(),
      .F2A_T_15_6(),
      .F2A_T_15_7(),
      .F2A_T_15_8(),
      .F2A_T_15_9(),
      .F2A_T_16_0(),
      .F2A_T_16_1(),
      .F2A_T_16_10(),
      .F2A_T_16_11(),
      .F2A_T_16_12(),
      .F2A_T_16_13(),
      .F2A_R_16_14(),
      .F2A_R_16_15(),
      .F2A_R_16_16(),
      .F2A_T_16_17(),
      .F2A_T_16_2(),
      .F2A_T_16_3(),
      .F2A_T_16_4(),
      .F2A_T_16_5(),
      .F2A_T_16_6(),
      .F2A_T_16_7(),
      .F2A_T_16_8(),
      .F2A_T_16_9(),
      .F2A_T_17_0(tcdm_clk_p2_int),
      .F2A_T_17_1(tcdm_req_p2),
      .F2A_T_17_10(tcdm_addr_p2[2]),
      .F2A_T_17_11(tcdm_addr_p2[3]),
      .F2A_T_17_2(tcdm_wen_p2),
      .F2A_T_17_3(tcdm_be_p2[0]),
      .F2A_T_17_4(tcdm_be_p2[1]),
      .F2A_T_17_5(tcdm_be_p2[2]),
      .F2A_T_17_6(tcdm_be_p2[3]),
      .F2A_T_17_7(),
      .F2A_T_17_8(tcdm_addr_p2[0]),
      .F2A_T_17_9(tcdm_addr_p2[1]),
      .F2A_T_18_0(tcdm_wdata_p2[0]),
      .F2A_T_18_1(tcdm_wdata_p2[1]),
      .F2A_T_18_10(tcdm_addr_p2[5]),
      .F2A_T_18_11(tcdm_addr_p2[6]),
      .F2A_T_18_12(tcdm_addr_p2[7]),
      .F2A_T_18_13(tcdm_addr_p2[8]),
      .F2A_T_18_14(tcdm_addr_p2[9]),
      .F2A_T_18_15(),
      .F2A_T_18_16(),
      .F2A_T_18_17(),
      .F2A_T_18_2(tcdm_wdata_p2[2]),
      .F2A_T_18_3(tcdm_wdata_p2[3]),
      .F2A_T_18_4(tcdm_wdata_p2[4]),
      .F2A_T_18_5(tcdm_wdata_p2[5]),
      .F2A_T_18_6(tcdm_wdata_p2[6]),
      .F2A_T_18_7(tcdm_wdata_p2[7]),
      .F2A_T_18_8(),
      .F2A_T_18_9(tcdm_addr_p2[4]),
      .F2A_T_19_0(tcdm_wdata_p2[8]),
      .F2A_T_19_1(tcdm_wdata_p2[9]),
      .F2A_T_19_10(tcdm_addr_p2[12]),
      .F2A_T_19_11(tcdm_addr_p2[13]),
      .F2A_T_19_2(tcdm_wdata_p2[10]),
      .F2A_T_19_3(tcdm_wdata_p2[11]),
      .F2A_T_19_4(tcdm_wdata_p2[12]),
      .F2A_T_19_5(tcdm_wdata_p2[13]),
      .F2A_T_19_6(tcdm_wdata_p2[14]),
      .F2A_T_19_7(tcdm_wdata_p2[15]),
      .F2A_T_19_8(tcdm_addr_p2[10]),
      .F2A_T_19_9(tcdm_addr_p2[11]),
      .F2A_T_1_0(),
      .F2A_T_1_1(),
      .F2A_T_1_10(),
      .F2A_T_1_11(),
      .F2A_T_1_2(),
      .F2A_T_1_3(),
      .F2A_T_1_4(),
      .F2A_T_1_5(),
      .F2A_T_1_6(),
      .F2A_T_1_7(),
      .F2A_T_1_8(),
      .F2A_T_1_9(),
      .F2A_T_20_0(tcdm_wdata_p2[16]),
      .F2A_T_20_1(tcdm_wdata_p2[17]),
      .F2A_T_20_10(),
      .F2A_T_20_11(),
      .F2A_T_20_12(tcdm_addr_p2[14]),
      .F2A_T_20_13(tcdm_addr_p2[15]),
      .F2A_T_20_14(tcdm_addr_p2[16]),
      .F2A_T_20_15(tcdm_addr_p2[17]),
      .F2A_T_20_16(tcdm_addr_p2[18]),
      .F2A_T_20_17(tcdm_addr_p2[19]),
      .F2A_T_20_2(tcdm_wdata_p2[18]),
      .F2A_T_20_3(tcdm_wdata_p2[19]),
      .F2A_T_20_4(tcdm_wdata_p2[20]),
      .F2A_T_20_5(tcdm_wdata_p2[21]),
      .F2A_T_20_6(tcdm_wdata_p2[22]),
      .F2A_T_20_7(tcdm_wdata_p2[23]),
      .F2A_T_20_8(),
      .F2A_T_20_9(),
      .F2A_T_21_0(tcdm_wdata_p2[24]),
      .F2A_T_21_1(tcdm_wdata_p2[25]),
      .F2A_T_21_10(),
      .F2A_T_21_11(),
      .F2A_T_21_2(tcdm_wdata_p2[26]),
      .F2A_T_21_3(tcdm_wdata_p2[27]),
      .F2A_T_21_4(tcdm_wdata_p2[28]),
      .F2A_T_21_5(tcdm_wdata_p2[29]),
      .F2A_T_21_6(tcdm_wdata_p2[30]),
      .F2A_T_21_7(tcdm_wdata_p2[31]),
      .F2A_T_21_8(),
      .F2A_T_21_9(),
      .F2A_T_22_0(),
      .F2A_T_22_1(),
      .F2A_T_22_10(),
      .F2A_T_22_11(),
      .F2A_T_22_12(),
      .F2A_T_22_13(),
      .F2A_T_22_14(),
      .F2A_T_22_15(),
      .F2A_T_22_16(),
      .F2A_T_22_17(),
      .F2A_T_22_2(),
      .F2A_T_22_3(),
      .F2A_T_22_4(),
      .F2A_T_22_5(),
      .F2A_T_22_6(),
      .F2A_T_22_7(),
      .F2A_T_22_8(),
      .F2A_T_22_9(),
      .F2A_T_23_0(tcdm_clk_p3_int),
      .F2A_T_23_1(tcdm_req_p3),
      .F2A_T_23_10(tcdm_addr_p3[2]),
      .F2A_T_23_11(tcdm_addr_p3[3]),
      .F2A_T_23_2(tcdm_wen_p3),
      .F2A_T_23_3(tcdm_be_p3[0]),
      .F2A_T_23_4(tcdm_be_p3[1]),
      .F2A_T_23_5(tcdm_be_p3[2]),
      .F2A_T_23_6(tcdm_be_p3[3]),
      .F2A_T_23_7(),
      .F2A_T_23_8(tcdm_addr_p3[0]),
      .F2A_T_23_9(tcdm_addr_p3[1]),
      .F2A_T_24_0(tcdm_wdata_p3[0]),
      .F2A_T_24_1(tcdm_wdata_p3[1]),
      .F2A_T_24_10(tcdm_addr_p3[5]),
      .F2A_T_24_11(tcdm_addr_p3[6]),
      .F2A_T_24_12(tcdm_addr_p3[7]),
      .F2A_T_24_13(tcdm_addr_p3[8]),
      .F2A_T_24_14(tcdm_addr_p3[9]),
      .F2A_T_24_15(),
      .F2A_T_24_16(),
      .F2A_T_24_17(),
      .F2A_T_24_2(tcdm_wdata_p3[2]),
      .F2A_T_24_3(tcdm_wdata_p3[3]),
      .F2A_T_24_4(tcdm_wdata_p3[4]),
      .F2A_T_24_5(tcdm_wdata_p3[5]),
      .F2A_T_24_6(tcdm_wdata_p3[6]),
      .F2A_T_24_7(tcdm_wdata_p3[7]),
      .F2A_T_24_8(),
      .F2A_T_24_9(tcdm_addr_p3[4]),
      .F2A_T_25_0(tcdm_wdata_p3[8]),
      .F2A_T_25_1(tcdm_wdata_p3[9]),
      .F2A_T_25_10(tcdm_addr_p3[12]),
      .F2A_T_25_11(tcdm_addr_p3[13]),
      .F2A_T_25_2(tcdm_wdata_p3[10]),
      .F2A_T_25_3(tcdm_wdata_p3[11]),
      .F2A_T_25_4(tcdm_wdata_p3[12]),
      .F2A_T_25_5(tcdm_wdata_p3[13]),
      .F2A_T_25_6(tcdm_wdata_p3[14]),
      .F2A_T_25_7(tcdm_wdata_p3[15]),
      .F2A_T_25_8(tcdm_addr_p3[10]),
      .F2A_T_25_9(tcdm_addr_p3[11]),
      .F2A_T_26_0(tcdm_wdata_p3[16]),
      .F2A_T_26_1(tcdm_wdata_p3[17]),
      .F2A_T_26_10(),
      .F2A_T_26_11(),
      .F2A_T_26_12(tcdm_addr_p3[14]),
      .F2A_T_26_13(tcdm_addr_p3[15]),
      .F2A_T_26_14(tcdm_addr_p3[16]),
      .F2A_T_26_15(tcdm_addr_p3[17]),
      .F2A_T_26_16(tcdm_addr_p3[18]),
      .F2A_T_26_17(tcdm_addr_p3[19]),
      .F2A_T_26_2(tcdm_wdata_p3[18]),
      .F2A_T_26_3(tcdm_wdata_p3[19]),
      .F2A_T_26_4(tcdm_wdata_p3[20]),
      .F2A_T_26_5(tcdm_wdata_p3[21]),
      .F2A_T_26_6(tcdm_wdata_p3[22]),
      .F2A_T_26_7(tcdm_wdata_p3[23]),
      .F2A_T_26_8(),
      .F2A_T_26_9(),
      .F2A_T_27_0(tcdm_wdata_p3[24]),
      .F2A_T_27_1(tcdm_wdata_p3[25]),
      .F2A_T_27_10(),
      .F2A_T_27_11(),
      .F2A_T_27_2(tcdm_wdata_p3[26]),
      .F2A_T_27_3(tcdm_wdata_p3[27]),
      .F2A_T_27_4(tcdm_wdata_p3[28]),
      .F2A_T_27_5(tcdm_wdata_p3[29]),
      .F2A_T_27_6(tcdm_wdata_p3[30]),
      .F2A_T_27_7(tcdm_wdata_p3[31]),
      .F2A_T_27_8(),
      .F2A_T_27_9(),
      .F2A_T_28_0(),
      .F2A_T_28_1(),
      .F2A_T_28_10(),
      .F2A_T_28_11(),
      .F2A_T_28_12(),
      .F2A_T_28_13(),
      .F2A_T_28_14(),
      .F2A_T_28_15(),
      .F2A_T_28_16(),
      .F2A_T_28_17(),
      .F2A_T_28_2(),
      .F2A_T_28_3(),
      .F2A_T_28_4(),
      .F2A_T_28_5(),
      .F2A_T_28_6(),
      .F2A_T_28_7(),
      .F2A_T_28_8(),
      .F2A_T_28_9(),
      .F2A_T_29_0(),
      .F2A_T_29_1(),
      .F2A_T_29_10(),
      .F2A_T_29_11(),
      .F2A_T_29_2(),
      .F2A_T_29_3(),
      .F2A_T_29_4(),
      .F2A_T_29_5(),
      .F2A_T_29_6(),
      .F2A_T_29_7(),
      .F2A_T_29_8(),
      .F2A_T_29_9(),
      .F2A_T_2_0(),
      .F2A_T_2_1(),
      .F2A_T_2_10(),
      .F2A_T_2_11(),
      .F2A_T_2_12(),
      .F2A_T_2_13(),
      .F2A_T_2_14(),
      .F2A_T_2_15(),
      .F2A_T_2_16(),
      .F2A_T_2_17(),
      .F2A_T_2_2(),
      .F2A_T_2_3(),
      .F2A_T_2_4(),
      .F2A_T_2_5(),
      .F2A_T_2_6(),
      .F2A_T_2_7(),
      .F2A_T_2_8(),
      .F2A_T_2_9(),
      .F2A_T_30_0(),
      .F2A_T_30_1(),
      .F2A_T_30_10(),
      .F2A_T_30_11(),
      .F2A_T_30_12(),
      .F2A_T_30_13(),
      .F2A_T_30_14(),
      .F2A_T_30_15(),
      .F2A_T_30_16(),
      .F2A_T_30_17(),
      .F2A_T_30_2(),
      .F2A_T_30_3(),
      .F2A_T_30_4(),
      .F2A_T_30_5(),
      .F2A_T_30_6(),
      .F2A_T_30_7(),
      .F2A_T_30_8(),
      .F2A_T_30_9(),
      .F2A_T_31_0(),
      .F2A_T_31_1(),
      .F2A_T_31_10(),
      .F2A_T_31_11(),
      .F2A_T_31_2(),
      .F2A_T_31_3(),
      .F2A_T_31_4(),
      .F2A_T_31_5(),
      .F2A_T_31_6(),
      .F2A_T_31_7(),
      .F2A_T_31_8(),
      .F2A_T_31_9(),
      .F2A_T_32_0(),
      .F2A_T_32_1(),
      .F2A_T_32_10(),
      .F2A_T_32_11(),
      .F2A_T_32_12(),
      .F2A_T_32_13(),
      .F2A_T_32_14(),
      .F2A_T_32_15(),
      .F2A_T_32_16(),
      .F2A_T_32_17(),
      .F2A_T_32_2(),
      .F2A_T_32_3(),
      .F2A_T_32_4(),
      .F2A_T_32_5(),
      .F2A_T_32_6(),
      .F2A_T_32_7(),
      .F2A_T_32_8(),
      .F2A_T_32_9(),
      .F2A_T_3_0(tcdm_clk_p0_int),
      .F2A_T_3_1(tcdm_req_p0),
      .F2A_T_3_10(tcdm_addr_p0[2]),
      .F2A_T_3_11(tcdm_addr_p0[3]),
      .F2A_T_3_2(tcdm_wen_p0),
      .F2A_T_3_3(tcdm_be_p0[0]),
      .F2A_T_3_4(tcdm_be_p0[1]),
      .F2A_T_3_5(tcdm_be_p0[2]),
      .F2A_T_3_6(tcdm_be_p0[3]),
      .F2A_T_3_7(),
      .F2A_T_3_8(tcdm_addr_p0[0]),
      .F2A_T_3_9(tcdm_addr_p0[1]),
      .F2A_T_4_0(tcdm_wdata_p0[0]),
      .F2A_T_4_1(tcdm_wdata_p0[1]),
      .F2A_T_4_10(tcdm_addr_p0[5]),
      .F2A_T_4_11(tcdm_addr_p0[6]),
      .F2A_T_4_12(tcdm_addr_p0[7]),
      .F2A_T_4_13(tcdm_addr_p0[8]),
      .F2A_T_4_14(tcdm_addr_p0[9]),
      .F2A_T_4_15(),
      .F2A_T_4_16(),
      .F2A_T_4_17(),
      .F2A_T_4_2(tcdm_wdata_p0[2]),
      .F2A_T_4_3(tcdm_wdata_p0[3]),
      .F2A_T_4_4(tcdm_wdata_p0[4]),
      .F2A_T_4_5(tcdm_wdata_p0[5]),
      .F2A_T_4_6(tcdm_wdata_p0[6]),
      .F2A_T_4_7(tcdm_wdata_p0[7]),
      .F2A_T_4_8(),
      .F2A_T_4_9(tcdm_addr_p0[4]),
      .F2A_T_5_0(tcdm_wdata_p0[8]),
      .F2A_T_5_1(tcdm_wdata_p0[9]),
      .F2A_T_5_10(tcdm_addr_p0[12]),
      .F2A_T_5_11(tcdm_addr_p0[13]),
      .F2A_T_5_2(tcdm_wdata_p0[10]),
      .F2A_T_5_3(tcdm_wdata_p0[11]),
      .F2A_T_5_4(tcdm_wdata_p0[12]),
      .F2A_T_5_5(tcdm_wdata_p0[13]),
      .F2A_T_5_6(tcdm_wdata_p0[14]),
      .F2A_T_5_7(tcdm_wdata_p0[15]),
      .F2A_T_5_8(tcdm_addr_p0[10]),
      .F2A_T_5_9(tcdm_addr_p0[11]),
      .F2A_T_6_0(tcdm_wdata_p0[16]),
      .F2A_T_6_1(tcdm_wdata_p0[17]),
      .F2A_T_6_10(),
      .F2A_T_6_11(),
      .F2A_T_6_12(tcdm_addr_p0[14]),
      .F2A_T_6_13(tcdm_addr_p0[15]),
      .F2A_T_6_14(tcdm_addr_p0[16]),
      .F2A_T_6_15(tcdm_addr_p0[17]),
      .F2A_T_6_16(tcdm_addr_p0[18]),
      .F2A_T_6_17(tcdm_addr_p0[19]),
      .F2A_T_6_2(tcdm_wdata_p0[18]),
      .F2A_T_6_3(tcdm_wdata_p0[19]),
      .F2A_T_6_4(tcdm_wdata_p0[20]),
      .F2A_T_6_5(tcdm_wdata_p0[21]),
      .F2A_T_6_6(tcdm_wdata_p0[22]),
      .F2A_T_6_7(tcdm_wdata_p0[23]),
      .F2A_T_6_8(),
      .F2A_T_6_9(),
      .F2A_T_7_0(tcdm_wdata_p0[24]),
      .F2A_T_7_1(tcdm_wdata_p0[25]),
      .F2A_T_7_10(),
      .F2A_T_7_11(),
      .F2A_T_7_2(tcdm_wdata_p0[26]),
      .F2A_T_7_3(tcdm_wdata_p0[27]),
      .F2A_T_7_4(tcdm_wdata_p0[28]),
      .F2A_T_7_5(tcdm_wdata_p0[29]),
      .F2A_T_7_6(tcdm_wdata_p0[30]),
      .F2A_T_7_7(tcdm_wdata_p0[31]),
      .F2A_T_7_8(),
      .F2A_T_7_9(),
      .F2A_T_8_0(),
      .F2A_T_8_1(),
      .F2A_T_8_10(),
      .F2A_T_8_11(),
      .F2A_T_8_12(),
      .F2A_T_8_13(),
      .F2A_T_8_14(),
      .F2A_T_8_15(),
      .F2A_T_8_16(),
      .F2A_T_8_17(),
      .F2A_T_8_2(),
      .F2A_T_8_3(),
      .F2A_T_8_4(),
      .F2A_T_8_5(),
      .F2A_T_8_6(),
      .F2A_T_8_7(),
      .F2A_T_8_8(),
      .F2A_T_8_9(),
      .F2A_T_9_0(tcdm_clk_p1_int),
      .F2A_T_9_1(tcdm_req_p1),
      .F2A_T_9_10(tcdm_addr_p1[2]),
      .F2A_T_9_11(tcdm_addr_p1[3]),
      .F2A_T_9_2(tcdm_wen_p1),
      .F2A_T_9_3(tcdm_be_p1[0]),
      .F2A_T_9_4(tcdm_be_p1[1]),
      .F2A_T_9_5(tcdm_be_p1[2]),
      .F2A_T_9_6(tcdm_be_p1[3]),
      .F2A_T_9_7(),
      .F2A_T_9_8(tcdm_addr_p1[0]),
      .F2A_T_9_9(tcdm_addr_p1[1]),
      .F2A_R_10_0(m0_m0_coef_in[20]),
      .F2A_R_10_1(m0_m0_coef_in[19]),
      .F2A_R_10_10(m0_m0_coef_in[10]),
      .F2A_R_10_11(m0_m0_coef_in[9]),
      .F2A_R_10_12(m0_m0_coef_in[8]),
      .F2A_R_10_13(m0_m0_coef_in[7]),
      .F2A_R_10_14(m0_m0_coef_in[6]),
      .F2A_R_10_15(m0_m0_coef_in[5]),
      .F2A_R_10_16(m0_m0_coef_in[4]),
      .F2A_R_10_17(m0_m0_coef_in[3]),
      .F2A_R_10_2(m0_m0_coef_in[18]),
      .F2A_R_10_3(m0_m0_coef_in[17]),
      .F2A_R_10_4(m0_m0_coef_in[16]),
      .F2A_R_10_5(m0_m0_coef_in[15]),
      .F2A_R_10_6(m0_m0_coef_in[14]),
      .F2A_R_10_7(m0_m0_coef_in[13]),
      .F2A_R_10_8(m0_m0_coef_in[12]),
      .F2A_R_10_9(m0_m0_coef_in[11]),
      .F2A_R_11_0(m0_m0_coef_in[2]),
      .F2A_R_11_1(m0_m0_coef_in[1]),
      .F2A_R_11_10(m0_coef_wdata[28]),
      .F2A_R_11_11(m0_coef_wdata[27]),
      .F2A_R_11_2(m0_m0_coef_in[0]),
      .F2A_R_11_3(m0_m0_mode[1]),
      .F2A_R_11_4(m0_m0_mode[0]),
      .F2A_R_11_5(m0_m0_tc),
      .F2A_R_11_6(m0_m0_reset),
      .F2A_R_11_7(m0_coef_wdata[31]),
      .F2A_R_11_8(m0_coef_wdata[30]),
      .F2A_R_11_9(m0_coef_wdata[29]),
      .F2A_R_12_0(m0_coef_wdata[26]),
      .F2A_R_12_1(m0_coef_wdata[25]),
      .F2A_R_12_10(m0_coef_wdata[16]),
      .F2A_R_12_11(m0_coef_wdata[15]),
      .F2A_R_12_12(m0_coef_wdata[14]),
      .F2A_R_12_13(m0_coef_wdata[13]),
      .F2A_R_12_14(m0_coef_wdata[12]),
      .F2A_R_12_15(m0_coef_wdata[11]),
      .F2A_R_12_16(m0_coef_wdata[10]),
      .F2A_R_12_17(m0_coef_wdata[9]),
      .F2A_R_12_2(m0_coef_wdata[24]),
      .F2A_R_12_3(m0_coef_wdata[23]),
      .F2A_R_12_4(m0_coef_wdata[22]),
      .F2A_R_12_5(m0_coef_wdata[21]),
      .F2A_R_12_6(m0_coef_wdata[20]),
      .F2A_R_12_7(m0_coef_wdata[19]),
      .F2A_R_12_8(m0_coef_wdata[18]),
      .F2A_R_12_9(m0_coef_wdata[17]),
      .F2A_R_13_0(m0_coef_wclk_int),
      .F2A_R_13_1(m0_coef_wdata[8]),
      .F2A_R_13_10(m0_coef_waddr[11]),
      .F2A_R_13_11(m0_coef_waddr[10]),
      .F2A_R_13_2(m0_coef_wdata[7]),
      .F2A_R_13_3(m0_coef_wdata[6]),
      .F2A_R_13_4(m0_coef_wdata[5]),
      .F2A_R_13_5(m0_coef_wdata[4]),
      .F2A_R_13_6(m0_coef_wdata[3]),
      .F2A_R_13_7(m0_coef_wdata[2]),
      .F2A_R_13_8(m0_coef_wdata[1]),
      .F2A_R_13_9(m0_coef_wdata[0]),
      .F2A_R_14_0(m0_coef_waddr[9]),
      .F2A_R_14_1(m0_coef_waddr[8]),
      .F2A_R_14_10(m0_coef_we),
      .F2A_R_14_11(m0_coef_wdsel),
      .F2A_R_14_12(m0_coef_rmode[1]),
      .F2A_R_14_13(m0_coef_rmode[0]),
      .F2A_R_14_14(m0_coef_raddr[11]),
      .F2A_R_14_15(m0_coef_raddr[10]),
      .F2A_R_14_16(m0_coef_raddr[9]),
      .F2A_R_14_17(m0_coef_raddr[8]),
      .F2A_R_14_2(m0_coef_waddr[7]),
      .F2A_R_14_3(m0_coef_waddr[6]),
      .F2A_R_14_4(m0_coef_waddr[5]),
      .F2A_R_14_5(m0_coef_waddr[4]),
      .F2A_R_14_6(m0_coef_waddr[3]),
      .F2A_R_14_7(m0_coef_waddr[2]),
      .F2A_R_14_8(m0_coef_waddr[1]),
      .F2A_R_14_9(m0_coef_waddr[0]),
      .F2A_R_15_0(m0_coef_rclk_int),
      .F2A_R_15_1(m0_coef_raddr[7]),
      .F2A_R_15_10(m0_coef_wmode[0]),
      .F2A_R_15_11(),
      .F2A_R_15_2(m0_coef_raddr[6]),
      .F2A_R_15_3(m0_coef_raddr[5]),
      .F2A_R_15_4(m0_coef_raddr[4]),
      .F2A_R_15_5(m0_coef_raddr[3]),
      .F2A_R_15_6(m0_coef_raddr[2]),
      .F2A_R_15_7(m0_coef_raddr[1]),
      .F2A_R_15_8(m0_coef_raddr[0]),
      .F2A_R_15_9(m0_coef_wmode[1]),
      .F2A_R_16_0(),
      .F2A_R_16_1(),
      .F2A_R_16_10(),
      .F2A_R_16_11(),
      .F2A_R_16_12(),
      .F2A_R_16_13(),
      .F2A_R_16_17(),
      .F2A_R_16_2(),
      .F2A_R_16_3(),
      .F2A_R_16_4(),
      .F2A_R_16_5(),
      .F2A_R_16_6(),
      .F2A_R_16_7(),
      .F2A_R_16_8(),
      .F2A_R_16_9(),
      .F2A_R_17_0(),
      .F2A_R_17_1(),
      .F2A_R_17_10(),
      .F2A_R_17_11(),
      .F2A_R_17_2(),
      .F2A_R_17_3(),
      .F2A_R_17_4(),
      .F2A_R_17_5(),
      .F2A_R_17_6(),
      .F2A_R_17_7(),
      .F2A_R_17_8(),
      .F2A_R_17_9(),
      .F2A_R_18_0(),
      .F2A_R_18_1(),
      .F2A_R_18_10(m0_m1_outsel[3]),
      .F2A_R_18_11(m0_m1_outsel[2]),
      .F2A_R_18_12(m0_m1_outsel[1]),
      .F2A_R_18_13(m0_m1_outsel[0]),
      .F2A_R_18_14(m0_m1_sat),
      .F2A_R_18_15(m0_m1_rnd),
      .F2A_R_18_16(m0_m1_clr),
      .F2A_R_18_17(m0_m1_clken),
      .F2A_R_18_2(),
      .F2A_R_18_3(),
      .F2A_R_18_4(),
      .F2A_R_18_5(),
      .F2A_R_18_6(),
      .F2A_R_18_7(),
      .F2A_R_18_8(m0_m1_outsel[5]),
      .F2A_R_18_9(m0_m1_outsel[4]),
      .F2A_R_19_0(m0_m1_clk_int),
      .F2A_R_19_1(m0_m1_osel),
      .F2A_R_19_10(m0_m1_coef_in[25]),
      .F2A_R_19_11(m0_m1_coef_in[24]),
      .F2A_R_19_2(m0_m1_tc),
      .F2A_R_19_3(m0_m1_reset),
      .F2A_R_19_4(m0_m1_coef_in[31]),
      .F2A_R_19_5(m0_m1_coef_in[30]),
      .F2A_R_19_6(m0_m1_coef_in[29]),
      .F2A_R_19_7(m0_m1_coef_in[28]),
      .F2A_R_19_8(m0_m1_coef_in[27]),
      .F2A_R_19_9(m0_m1_coef_in[26]),
      .F2A_R_1_0(),
      .F2A_R_1_1(),
      .F2A_R_1_10(),
      .F2A_R_1_11(),
      .F2A_R_1_2(),
      .F2A_R_1_3(),
      .F2A_R_1_4(),
      .F2A_R_1_5(),
      .F2A_R_1_6(),
      .F2A_R_1_7(),
      .F2A_R_1_8(),
      .F2A_R_1_9(),
      .F2A_R_20_0(m0_m1_coef_in[23]),
      .F2A_R_20_1(m0_m1_coef_in[22]),
      .F2A_R_20_10(m0_m1_coef_in[13]),
      .F2A_R_20_11(m0_m1_coef_in[12]),
      .F2A_R_20_12(m0_m1_coef_in[11]),
      .F2A_R_20_13(m0_m1_coef_in[10]),
      .F2A_R_20_14(m0_m1_coef_in[9]),
      .F2A_R_20_15(m0_m1_coef_in[8]),
      .F2A_R_20_16(m0_m1_coef_in[7]),
      .F2A_R_20_17(m0_m1_coef_in[6]),
      .F2A_R_20_2(m0_m1_coef_in[21]),
      .F2A_R_20_3(m0_m1_coef_in[20]),
      .F2A_R_20_4(m0_m1_coef_in[19]),
      .F2A_R_20_5(m0_m1_coef_in[18]),
      .F2A_R_20_6(m0_m1_coef_in[17]),
      .F2A_R_20_7(m0_m1_coef_in[16]),
      .F2A_R_20_8(m0_m1_coef_in[15]),
      .F2A_R_20_9(m0_m1_coef_in[14]),
      .F2A_R_21_0(m0_m1_coef_in[5]),
      .F2A_R_21_1(m0_m1_coef_in[4]),
      .F2A_R_21_10(m0_m1_oper_in[30]),
      .F2A_R_21_11(m0_m1_oper_in[29]),
      .F2A_R_21_2(m0_m1_coef_in[3]),
      .F2A_R_21_3(m0_m1_coef_in[2]),
      .F2A_R_21_4(m0_m1_coef_in[1]),
      .F2A_R_21_5(m0_m1_coef_in[0]),
      .F2A_R_21_6(m0_m1_mode[1]),
      .F2A_R_21_7(m0_m1_csel),
      .F2A_R_21_8(m0_m1_mode[0]),
      .F2A_R_21_9(m0_m1_oper_in[31]),
      .F2A_R_22_0(m0_m1_oper_in[28]),
      .F2A_R_22_1(m0_m1_oper_in[27]),
      .F2A_R_22_10(m0_m1_oper_in[18]),
      .F2A_R_22_11(m0_m1_oper_in[17]),
      .F2A_R_22_12(m0_m1_oper_in[16]),
      .F2A_R_22_13(m0_m1_oper_in[15]),
      .F2A_R_22_14(m0_m1_oper_in[14]),
      .F2A_R_22_15(m0_m1_oper_in[13]),
      .F2A_R_22_16(m0_m1_oper_in[12]),
      .F2A_R_22_17(m0_m1_oper_in[11]),
      .F2A_R_22_2(m0_m1_oper_in[26]),
      .F2A_R_22_3(m0_m1_oper_in[25]),
      .F2A_R_22_4(m0_m1_oper_in[24]),
      .F2A_R_22_5(m0_m1_oper_in[23]),
      .F2A_R_22_6(m0_m1_oper_in[22]),
      .F2A_R_22_7(m0_m1_oper_in[21]),
      .F2A_R_22_8(m0_m1_oper_in[20]),
      .F2A_R_22_9(m0_m1_oper_in[19]),
      .F2A_R_23_0(m0_m1_oper_in[10]),
      .F2A_R_23_1(m0_m1_oper_in[9]),
      .F2A_R_23_10(m0_m1_oper_in[0]),
      .F2A_R_23_11(),
      .F2A_R_23_2(m0_m1_oper_in[8]),
      .F2A_R_23_3(m0_m1_oper_in[7]),
      .F2A_R_23_4(m0_m1_oper_in[6]),
      .F2A_R_23_5(m0_m1_oper_in[5]),
      .F2A_R_23_6(m0_m1_oper_in[4]),
      .F2A_R_23_7(m0_m1_oper_in[3]),
      .F2A_R_23_8(m0_m1_oper_in[2]),
      .F2A_R_23_9(m0_m1_oper_in[1]),
      .F2A_R_24_0(),
      .F2A_R_24_1(),
      .F2A_R_24_10(),
      .F2A_R_24_11(),
      .F2A_R_24_12(),
      .F2A_R_24_13(),
      .F2A_R_24_14(),
      .F2A_R_24_15(),
      .F2A_R_24_16(m0_oper1_wdata[31]),
      .F2A_R_24_17(m0_oper1_wdata[30]),
      .F2A_R_24_2(),
      .F2A_R_24_3(),
      .F2A_R_24_4(),
      .F2A_R_24_5(),
      .F2A_R_24_6(),
      .F2A_R_24_7(),
      .F2A_R_24_8(),
      .F2A_R_24_9(),
      .F2A_R_25_0(m0_oper1_wdata[29]),
      .F2A_R_25_1(m0_oper1_wdata[28]),
      .F2A_R_25_10(m0_oper1_wdata[19]),
      .F2A_R_25_11(m0_oper1_wdata[18]),
      .F2A_R_25_2(m0_oper1_wdata[27]),
      .F2A_R_25_3(m0_oper1_wdata[26]),
      .F2A_R_25_4(m0_oper1_wdata[25]),
      .F2A_R_25_5(m0_oper1_wdata[24]),
      .F2A_R_25_6(m0_oper1_wdata[23]),
      .F2A_R_25_7(m0_oper1_wdata[22]),
      .F2A_R_25_8(m0_oper1_wdata[21]),
      .F2A_R_25_9(m0_oper1_wdata[20]),
      .F2A_R_26_0(m0_oper1_wdata[17]),
      .F2A_R_26_1(m0_oper1_wdata[16]),
      .F2A_R_26_10(m0_oper1_wdata[7]),
      .F2A_R_26_11(m0_oper1_wdata[6]),
      .F2A_R_26_12(m0_oper1_wdata[5]),
      .F2A_R_26_13(m0_oper1_wdata[4]),
      .F2A_R_26_14(m0_oper1_wdata[3]),
      .F2A_R_26_15(m0_oper1_wdata[2]),
      .F2A_R_26_16(m0_oper1_wdata[1]),
      .F2A_R_26_17(m0_oper1_wdata[0]),
      .F2A_R_26_2(m0_oper1_wdata[15]),
      .F2A_R_26_3(m0_oper1_wdata[14]),
      .F2A_R_26_4(m0_oper1_wdata[13]),
      .F2A_R_26_5(m0_oper1_wdata[12]),
      .F2A_R_26_6(m0_oper1_wdata[11]),
      .F2A_R_26_7(m0_oper1_wdata[10]),
      .F2A_R_26_8(m0_oper1_wdata[9]),
      .F2A_R_26_9(m0_oper1_wdata[8]),
      .F2A_R_27_0(m0_oper1_waddr[11]),
      .F2A_R_27_1(m0_oper1_waddr[10]),
      .F2A_R_27_10(m0_oper1_waddr[1]),
      .F2A_R_27_11(m0_oper1_waddr[0]),
      .F2A_R_27_2(m0_oper1_waddr[9]),
      .F2A_R_27_3(m0_oper1_waddr[8]),
      .F2A_R_27_4(m0_oper1_waddr[7]),
      .F2A_R_27_5(m0_oper1_waddr[6]),
      .F2A_R_27_6(m0_oper1_waddr[5]),
      .F2A_R_27_7(m0_oper1_waddr[4]),
      .F2A_R_27_8(m0_oper1_waddr[3]),
      .F2A_R_27_9(m0_oper1_waddr[2]),
      .F2A_R_28_0(m0_oper1_wclk_int),
      .F2A_R_28_1(m0_oper1_wmode[1]),
      .F2A_R_28_10(),
      .F2A_R_28_11(),
      .F2A_R_28_12(),
      .F2A_R_28_13(),
      .F2A_R_28_14(),
      .F2A_R_28_15(m0_oper1_rmode[1]),
      .F2A_R_28_16(m0_oper1_rmode[0]),
      .F2A_R_28_17(m0_oper1_raddr[11]),
      .F2A_R_28_2(m0_oper1_wmode[0]),
      .F2A_R_28_3(m0_oper1_wdsel),
      .F2A_R_28_4(m0_oper1_we),
      .F2A_R_28_5(),
      .F2A_R_28_6(),
      .F2A_R_28_7(),
      .F2A_R_28_8(),
      .F2A_R_28_9(),
      .F2A_R_29_0(m0_oper1_rclk_int),
      .F2A_R_29_1(m0_oper1_raddr[10]),
      .F2A_R_29_10(m0_oper1_raddr[1]),
      .F2A_R_29_11(m0_oper1_raddr[0]),
      .F2A_R_29_2(m0_oper1_raddr[9]),
      .F2A_R_29_3(m0_oper1_raddr[8]),
      .F2A_R_29_4(m0_oper1_raddr[7]),
      .F2A_R_29_5(m0_oper1_raddr[6]),
      .F2A_R_29_6(m0_oper1_raddr[5]),
      .F2A_R_29_7(m0_oper1_raddr[4]),
      .F2A_R_29_8(m0_oper1_raddr[3]),
      .F2A_R_29_9(m0_oper1_raddr[2]),
      .F2A_R_2_0(m0_oper0_wclk_int),
      .F2A_R_2_1(m0_oper0_wmode[1]),
      .F2A_R_2_10(m0_oper0_wdata[27]),
      .F2A_R_2_11(m0_oper0_wdata[26]),
      .F2A_R_2_12(m0_oper0_wdata[25]),
      .F2A_R_2_13(m0_oper0_wdata[24]),
      .F2A_R_2_14(m0_oper0_wdata[23]),
      .F2A_R_2_15(m0_oper0_wdata[22]),
      .F2A_R_2_16(m0_oper0_wdata[21]),
      .F2A_R_2_17(m0_oper0_wdata[20]),
      .F2A_R_2_2(m0_oper0_wmode[0]),
      .F2A_R_2_3(m0_oper0_wdsel),
      .F2A_R_2_4(m0_oper0_rmode[1]),
      .F2A_R_2_5(m0_oper0_rmode[0]),
      .F2A_R_2_6(m0_oper0_wdata[31]),
      .F2A_R_2_7(m0_oper0_wdata[30]),
      .F2A_R_2_8(m0_oper0_wdata[29]),
      .F2A_R_2_9(m0_oper0_wdata[28]),
      .F2A_R_30_0(),
      .F2A_R_30_1(),
      .F2A_R_30_10(),
      .F2A_R_30_11(),
      .F2A_R_30_12(),
      .F2A_R_30_13(),
      .F2A_R_30_14(),
      .F2A_R_30_15(),
      .F2A_R_30_16(),
      .F2A_R_30_17(),
      .F2A_R_30_2(),
      .F2A_R_30_3(),
      .F2A_R_30_4(),
      .F2A_R_30_5(),
      .F2A_R_30_6(),
      .F2A_R_30_7(),
      .F2A_R_30_8(),
      .F2A_R_30_9(),
      .F2A_R_31_0(),
      .F2A_R_31_1(),
      .F2A_R_31_10(),
      .F2A_R_31_11(),
      .F2A_R_31_2(),
      .F2A_R_31_3(),
      .F2A_R_31_4(),
      .F2A_R_31_5(),
      .F2A_R_31_6(),
      .F2A_R_31_7(),
      .F2A_R_31_8(),
      .F2A_R_31_9(),
      .F2A_R_32_0(),
      .F2A_R_32_1(),
      .F2A_R_32_10(),
      .F2A_R_32_11(),
      .F2A_R_32_12(),
      .F2A_R_32_13(),
      .F2A_R_32_14(),
      .F2A_R_32_15(),
      .F2A_R_32_16(),
      .F2A_R_32_17(),
      .F2A_R_32_2(),
      .F2A_R_32_3(),
      .F2A_R_32_4(),
      .F2A_R_32_5(),
      .F2A_R_32_6(),
      .F2A_R_32_7(),
      .F2A_R_32_8(),
      .F2A_R_32_9(),
      .F2A_R_3_0(m0_oper0_wdata[19]),
      .F2A_R_3_1(m0_oper0_wdata[18]),
      .F2A_R_3_10(m0_oper0_wdata[9]),
      .F2A_R_3_11(m0_oper0_wdata[8]),
      .F2A_R_3_2(m0_oper0_wdata[17]),
      .F2A_R_3_3(m0_oper0_wdata[16]),
      .F2A_R_3_4(m0_oper0_wdata[15]),
      .F2A_R_3_5(m0_oper0_wdata[14]),
      .F2A_R_3_6(m0_oper0_wdata[13]),
      .F2A_R_3_7(m0_oper0_wdata[12]),
      .F2A_R_3_8(m0_oper0_wdata[11]),
      .F2A_R_3_9(m0_oper0_wdata[10]),
      .F2A_R_4_0(m0_oper0_wdata[7]),
      .F2A_R_4_1(m0_oper0_wdata[6]),
      .F2A_R_4_10(m0_oper0_waddr[9]),
      .F2A_R_4_11(m0_oper0_waddr[8]),
      .F2A_R_4_12(m0_oper0_waddr[7]),
      .F2A_R_4_13(m0_oper0_waddr[6]),
      .F2A_R_4_14(m0_oper0_waddr[5]),
      .F2A_R_4_15(m0_oper0_waddr[4]),
      .F2A_R_4_16(m0_oper0_waddr[3]),
      .F2A_R_4_17(m0_oper0_waddr[2]),
      .F2A_R_4_2(m0_oper0_wdata[5]),
      .F2A_R_4_3(m0_oper0_wdata[4]),
      .F2A_R_4_4(m0_oper0_wdata[3]),
      .F2A_R_4_5(m0_oper0_wdata[2]),
      .F2A_R_4_6(m0_oper0_wdata[1]),
      .F2A_R_4_7(m0_oper0_wdata[0]),
      .F2A_R_4_8(m0_oper0_waddr[11]),
      .F2A_R_4_9(m0_oper0_waddr[10]),
      .F2A_R_5_0(m0_oper0_waddr[1]),
      .F2A_R_5_1(m0_oper0_waddr[0]),
      .F2A_R_5_10(m0_oper0_raddr[4]),
      .F2A_R_5_11(m0_oper0_raddr[3]),
      .F2A_R_5_2(m0_oper0_we),
      .F2A_R_5_3(m0_oper0_raddr[11]),
      .F2A_R_5_4(m0_oper0_raddr[10]),
      .F2A_R_5_5(m0_oper0_raddr[9]),
      .F2A_R_5_6(m0_oper0_raddr[8]),
      .F2A_R_5_7(m0_oper0_raddr[7]),
      .F2A_R_5_8(m0_oper0_raddr[6]),
      .F2A_R_5_9(m0_oper0_raddr[5]),
      .F2A_R_6_0(m0_oper0_rclk_int),
      .F2A_R_6_1(m0_oper0_raddr[2]),
      .F2A_R_6_10(m0_m0_outsel[1]),
      .F2A_R_6_11(m0_m0_outsel[0]),
      .F2A_R_6_12(m0_m0_sat),
      .F2A_R_6_13(m0_m0_rnd),
      .F2A_R_6_14(m0_m0_clr),
      .F2A_R_6_15(m0_m0_oper_in[31]),
      .F2A_R_6_16(m0_m0_oper_in[30]),
      .F2A_R_6_17(m0_m0_oper_in[29]),
      .F2A_R_6_2(m0_oper0_raddr[1]),
      .F2A_R_6_3(m0_oper0_raddr[0]),
      .F2A_R_6_4(m0_m0_osel),
      .F2A_R_6_5(m0_m0_clken),
      .F2A_R_6_6(m0_m0_outsel[5]),
      .F2A_R_6_7(m0_m0_outsel[4]),
      .F2A_R_6_8(m0_m0_outsel[3]),
      .F2A_R_6_9(m0_m0_outsel[2]),
      .F2A_R_7_0(m0_m0_clk_int),
      .F2A_R_7_1(m0_m0_oper_in[28]),
      .F2A_R_7_10(m0_m0_oper_in[19]),
      .F2A_R_7_11(m0_m0_oper_in[18]),
      .F2A_R_7_2(m0_m0_oper_in[27]),
      .F2A_R_7_3(m0_m0_oper_in[26]),
      .F2A_R_7_4(m0_m0_oper_in[25]),
      .F2A_R_7_5(m0_m0_oper_in[24]),
      .F2A_R_7_6(m0_m0_oper_in[23]),
      .F2A_R_7_7(m0_m0_oper_in[22]),
      .F2A_R_7_8(m0_m0_oper_in[21]),
      .F2A_R_7_9(m0_m0_oper_in[20]),
      .F2A_R_8_0(m0_m0_oper_in[17]),
      .F2A_R_8_1(m0_m0_oper_in[16]),
      .F2A_R_8_10(m0_m0_oper_in[7]),
      .F2A_R_8_11(m0_m0_oper_in[6]),
      .F2A_R_8_12(m0_m0_oper_in[5]),
      .F2A_R_8_13(m0_m0_oper_in[4]),
      .F2A_R_8_14(m0_m0_oper_in[3]),
      .F2A_R_8_15(m0_m0_oper_in[2]),
      .F2A_R_8_16(m0_m0_oper_in[1]),
      .F2A_R_8_17(m0_m0_oper_in[0]),
      .F2A_R_8_2(m0_m0_oper_in[15]),
      .F2A_R_8_3(m0_m0_oper_in[14]),
      .F2A_R_8_4(m0_m0_oper_in[13]),
      .F2A_R_8_5(m0_m0_oper_in[12]),
      .F2A_R_8_6(m0_m0_oper_in[11]),
      .F2A_R_8_7(m0_m0_oper_in[10]),
      .F2A_R_8_8(m0_m0_oper_in[9]),
      .F2A_R_8_9(m0_m0_oper_in[8]),
      .F2A_R_9_0(m0_m0_csel),
      .F2A_R_9_1(m0_m0_coef_in[31]),
      .F2A_R_9_10(m0_m0_coef_in[22]),
      .F2A_R_9_11(m0_m0_coef_in[21]),
      .F2A_R_9_2(m0_m0_coef_in[30]),
      .F2A_R_9_3(m0_m0_coef_in[29]),
      .F2A_R_9_4(m0_m0_coef_in[28]),
      .F2A_R_9_5(m0_m0_coef_in[27]),
      .F2A_R_9_6(m0_m0_coef_in[26]),
      .F2A_R_9_7(m0_m0_coef_in[25]),
      .F2A_R_9_8(m0_m0_coef_in[24]),
      .F2A_R_9_9(m0_m0_coef_in[23]),
      .F2Adef_B_10_0(),
      .F2Adef_B_10_1(),
      .F2Adef_B_10_2(),
      .F2Adef_B_10_3(),
      .F2Adef_B_10_4(),
      .F2Adef_B_10_5(),
      .F2Adef_B_10_6(),
      .F2Adef_B_11_0(),
      .F2Adef_B_11_1(),
      .F2Adef_B_11_2(),
      .F2Adef_B_11_3(),
      .F2Adef_B_12_0(),
      .F2Adef_B_12_1(),
      .F2Adef_B_12_2(),
      .F2Adef_B_12_3(),
      .F2Adef_B_12_4(),
      .F2Adef_B_12_5(),
      .F2Adef_B_12_6(),
      .F2Adef_B_13_0(m1_coef_powerdn),
      .F2Adef_B_13_1(m1_coef_wclk_def),
      .F2Adef_B_13_2(),
      .F2Adef_B_13_3(),
      .F2Adef_B_14_0(),
      .F2Adef_B_14_1(),
      .F2Adef_B_14_2(),
      .F2Adef_B_14_3(),
      .F2Adef_B_14_4(),
      .F2Adef_B_14_5(),
      .F2Adef_B_14_6(),
      .F2Adef_B_15_0(m1_coef_rclk_def),
      .F2Adef_B_15_1(),
      .F2Adef_B_15_2(),
      .F2Adef_B_15_3(),
      .F2Adef_B_16_0(),
      .F2Adef_B_16_1(),
      .F2Adef_B_16_2(),
      .F2Adef_B_16_3(),
      .F2Adef_B_16_4(),
      .F2Adef_B_16_5(),
      .F2Adef_B_16_6(),
      .F2Adef_B_17_0(),
      .F2Adef_B_17_1(),
      .F2Adef_B_17_2(),
      .F2Adef_B_17_3(),
      .F2Adef_B_18_0(),
      .F2Adef_B_18_1(),
      .F2Adef_B_18_2(),
      .F2Adef_B_18_3(),
      .F2Adef_B_18_4(),
      .F2Adef_B_18_5(),
      .F2Adef_B_18_6(),
      .F2Adef_B_19_0(m1_m1_clk_def),
      .F2Adef_B_19_1(),
      .F2Adef_B_19_2(),
      .F2Adef_B_19_3(),
      .F2Adef_B_1_0(),
      .F2Adef_B_1_1(),
      .F2Adef_B_1_2(),
      .F2Adef_B_1_3(),
      .F2Adef_B_20_0(),
      .F2Adef_B_20_1(),
      .F2Adef_B_20_2(),
      .F2Adef_B_20_3(),
      .F2Adef_B_20_4(),
      .F2Adef_B_20_5(),
      .F2Adef_B_20_6(),
      .F2Adef_B_21_0(),
      .F2Adef_B_21_1(),
      .F2Adef_B_21_2(),
      .F2Adef_B_21_3(),
      .F2Adef_B_22_0(),
      .F2Adef_B_22_1(),
      .F2Adef_B_22_2(),
      .F2Adef_B_22_3(),
      .F2Adef_B_22_4(),
      .F2Adef_B_22_5(),
      .F2Adef_B_22_6(),
      .F2Adef_B_23_0(),
      .F2Adef_B_23_1(),
      .F2Adef_B_23_2(),
      .F2Adef_B_23_3(),
      .F2Adef_B_24_0(),
      .F2Adef_B_24_1(m1_oper1_powerdn),
      .F2Adef_B_24_2(),
      .F2Adef_B_24_3(),
      .F2Adef_B_24_4(),
      .F2Adef_B_24_5(),
      .F2Adef_B_24_6(),
      .F2Adef_B_25_0(),
      .F2Adef_B_25_1(),
      .F2Adef_B_25_2(),
      .F2Adef_B_25_3(),
      .F2Adef_B_26_0(),
      .F2Adef_B_26_1(),
      .F2Adef_B_26_2(),
      .F2Adef_B_26_3(),
      .F2Adef_B_26_4(),
      .F2Adef_B_26_5(),
      .F2Adef_B_26_6(),
      .F2Adef_B_27_0(),
      .F2Adef_B_27_1(),
      .F2Adef_B_27_2(),
      .F2Adef_B_27_3(),
      .F2Adef_B_28_0(m1_oper1_wclk_def),
      .F2Adef_B_28_1(),
      .F2Adef_B_28_2(),
      .F2Adef_B_28_3(),
      .F2Adef_B_28_4(),
      .F2Adef_B_28_5(),
      .F2Adef_B_28_6(),
      .F2Adef_B_29_0(m1_oper1_rclk_def),
      .F2Adef_B_29_1(),
      .F2Adef_B_29_2(),
      .F2Adef_B_29_3(),
      .F2Adef_B_2_0(m1_oper0_wclk_def),
      .F2Adef_B_2_1(),
      .F2Adef_B_2_2(),
      .F2Adef_B_2_3(),
      .F2Adef_B_2_4(),
      .F2Adef_B_2_5(),
      .F2Adef_B_2_6(),
      .F2Adef_B_30_0(),
      .F2Adef_B_30_1(),
      .F2Adef_B_30_2(),
      .F2Adef_B_30_3(),
      .F2Adef_B_30_4(),
      .F2Adef_B_30_5(),
      .F2Adef_B_30_6(),
      .F2Adef_B_31_0(),
      .F2Adef_B_31_1(),
      .F2Adef_B_31_2(),
      .F2Adef_B_31_3(),
      .F2Adef_B_32_0(),
      .F2Adef_B_32_1(),
      .F2Adef_B_32_2(),
      .F2Adef_B_32_3(),
      .F2Adef_B_32_4(),
      .F2Adef_B_32_5(),
      .F2Adef_B_32_6(),
      .F2Adef_B_3_0(),
      .F2Adef_B_3_1(),
      .F2Adef_B_3_2(),
      .F2Adef_B_3_3(),
      .F2Adef_B_4_0(),
      .F2Adef_B_4_1(),
      .F2Adef_B_4_2(),
      .F2Adef_B_4_3(),
      .F2Adef_B_4_4(),
      .F2Adef_B_4_5(),
      .F2Adef_B_4_6(),
      .F2Adef_B_5_0(),
      .F2Adef_B_5_1(),
      .F2Adef_B_5_2(),
      .F2Adef_B_5_3(),
      .F2Adef_B_6_0(m1_oper0_rclk_def),
      .F2Adef_B_6_1(m1_oper0_powerdn),
      .F2Adef_B_6_2(),
      .F2Adef_B_6_3(),
      .F2Adef_B_6_4(),
      .F2Adef_B_6_5(),
      .F2Adef_B_6_6(),
      .F2Adef_B_7_0(m1_m0_clk_def),
      .F2Adef_B_7_1(),
      .F2Adef_B_7_2(),
      .F2Adef_B_7_3(),
      .F2Adef_B_8_0(),
      .F2Adef_B_8_1(),
      .F2Adef_B_8_2(),
      .F2Adef_B_8_3(),
      .F2Adef_B_8_4(),
      .F2Adef_B_8_5(),
      .F2Adef_B_8_6(),
      .F2Adef_B_9_0(),
      .F2Adef_B_9_1(),
      .F2Adef_B_9_2(),
      .F2Adef_B_9_3(),
      .F2Adef_L_10_0(),
      .F2Adef_L_10_1(),
      .F2Adef_L_10_2(),
      .F2Adef_L_10_3(),
      .F2Adef_L_10_4(),
      .F2Adef_L_10_5(),
      .F2Adef_L_10_6(),
      .F2Adef_L_11_0(),
      .F2Adef_L_11_1(),
      .F2Adef_L_11_2(),
      .F2Adef_L_11_3(),
      .F2Adef_L_12_0(),
      .F2Adef_L_12_1(),
      .F2Adef_L_12_2(),
      .F2Adef_L_12_3(),
      .F2Adef_L_12_4(),
      .F2Adef_L_12_5(),
      .F2Adef_L_12_6(),
      .F2Adef_L_13_0(lint_clk_def),
      .F2Adef_L_13_1(),
      .F2Adef_L_13_2(),
      .F2Adef_L_13_3(),
      .F2Adef_L_14_0(),
      .F2Adef_L_14_1(),
      .F2Adef_L_14_2(),
      .F2Adef_L_14_3(),
      .F2Adef_L_14_4(),
      .F2Adef_L_14_5(),
      .F2Adef_L_14_6(),
      .F2Adef_L_15_0(),
      .F2Adef_L_15_1(),
      .F2Adef_L_15_2(),
      .F2Adef_L_15_3(),
      .F2Adef_L_16_0(),
      .F2Adef_L_16_1(),
      .F2Adef_L_16_2(),
      .F2Adef_L_16_3(),
      .F2Adef_L_16_4(),
      .F2Adef_L_16_5(),
      .F2Adef_L_16_6(),
      .F2Adef_L_17_0(),
      .F2Adef_L_17_1(),
      .F2Adef_L_17_2(),
      .F2Adef_L_17_3(),
      .F2Adef_L_18_0(),
      .F2Adef_L_18_1(),
      .F2Adef_L_18_2(),
      .F2Adef_L_18_3(),
      .F2Adef_L_18_4(),
      .F2Adef_L_18_5(),
      .F2Adef_L_18_6(),
      .F2Adef_L_19_0(),
      .F2Adef_L_19_1(),
      .F2Adef_L_19_2(),
      .F2Adef_L_19_3(),
      .F2Adef_L_1_0(),
      .F2Adef_L_1_1(),
      .F2Adef_L_1_2(),
      .F2Adef_L_1_3(),
      .F2Adef_L_20_0(),
      .F2Adef_L_20_1(),
      .F2Adef_L_20_2(),
      .F2Adef_L_20_3(),
      .F2Adef_L_20_4(),
      .F2Adef_L_20_5(),
      .F2Adef_L_20_6(),
      .F2Adef_L_21_0(),
      .F2Adef_L_21_1(),
      .F2Adef_L_21_2(),
      .F2Adef_L_21_3(),
      .F2Adef_L_22_0(),
      .F2Adef_L_22_1(),
      .F2Adef_L_22_2(),
      .F2Adef_L_22_3(),
      .F2Adef_L_22_4(),
      .F2Adef_L_22_5(),
      .F2Adef_L_22_6(),
      .F2Adef_L_23_0(),
      .F2Adef_L_23_1(),
      .F2Adef_L_23_2(),
      .F2Adef_L_23_3(),
      .F2Adef_L_24_0(),
      .F2Adef_L_24_1(),
      .F2Adef_L_24_2(),
      .F2Adef_L_24_3(),
      .F2Adef_L_24_4(),
      .F2Adef_L_24_5(),
      .F2Adef_L_24_6(),
      .F2Adef_L_25_0(),
      .F2Adef_L_25_1(),
      .F2Adef_L_25_2(),
      .F2Adef_L_25_3(),
      .F2Adef_L_26_0(),
      .F2Adef_L_26_1(),
      .F2Adef_L_26_2(),
      .F2Adef_L_26_3(),
      .F2Adef_L_26_4(),
      .F2Adef_L_26_5(),
      .F2Adef_L_26_6(),
      .F2Adef_L_27_0(),
      .F2Adef_L_27_1(),
      .F2Adef_L_27_2(),
      .F2Adef_L_27_3(),
      .F2Adef_L_28_0(),
      .F2Adef_L_28_1(),
      .F2Adef_L_28_2(),
      .F2Adef_L_28_3(),
      .F2Adef_L_28_4(),
      .F2Adef_L_28_5(),
      .F2Adef_L_28_6(),
      .F2Adef_L_29_0(),
      .F2Adef_L_29_1(),
      .F2Adef_L_29_2(),
      .F2Adef_L_29_3(),
      .F2Adef_L_2_0(version[0]),
      .F2Adef_L_2_1(version[1]),
      .F2Adef_L_2_2(version[2]),
      .F2Adef_L_2_3(version[3]),
      .F2Adef_L_2_4(version[4]),
      .F2Adef_L_2_5(version[5]),
      .F2Adef_L_2_6(version[6]),
      .F2Adef_L_30_0(),
      .F2Adef_L_30_1(),
      .F2Adef_L_30_2(),
      .F2Adef_L_30_3(),
      .F2Adef_L_30_4(),
      .F2Adef_L_30_5(),
      .F2Adef_L_30_6(),
      .F2Adef_L_31_0(),
      .F2Adef_L_31_1(),
      .F2Adef_L_31_2(),
      .F2Adef_L_31_3(),
      .F2Adef_L_32_0(),
      .F2Adef_L_32_1(),
      .F2Adef_L_32_2(),
      .F2Adef_L_32_3(),
      .F2Adef_L_32_4(),
      .F2Adef_L_32_5(),
      .F2Adef_L_32_6(),
      .F2Adef_L_3_0(),
      .F2Adef_L_3_1(),
      .F2Adef_L_3_2(),
      .F2Adef_L_3_3(),
      .F2Adef_L_4_0(version[7]),
      .F2Adef_L_4_1(),
      .F2Adef_L_4_2(),
      .F2Adef_L_4_3(),
      .F2Adef_L_4_4(),
      .F2Adef_L_4_5(),
      .F2Adef_L_4_6(),
      .F2Adef_L_5_0(),
      .F2Adef_L_5_1(),
      .F2Adef_L_5_2(),
      .F2Adef_L_5_3(),
      .F2Adef_L_6_0(),
      .F2Adef_L_6_1(),
      .F2Adef_L_6_2(),
      .F2Adef_L_6_3(),
      .F2Adef_L_6_4(),
      .F2Adef_L_6_5(),
      .F2Adef_L_6_6(),
      .F2Adef_L_7_0(),
      .F2Adef_L_7_1(),
      .F2Adef_L_7_2(),
      .F2Adef_L_7_3(),
      .F2Adef_L_8_0(),
      .F2Adef_L_8_1(),
      .F2Adef_L_8_2(),
      .F2Adef_L_8_3(),
      .F2Adef_L_8_4(),
      .F2Adef_L_8_5(),
      .F2Adef_L_8_6(),
      .F2Adef_L_9_0(),
      .F2Adef_L_9_1(),
      .F2Adef_L_9_2(),
      .F2Adef_L_9_3(),
      .F2Adef_T_10_0(),
      .F2Adef_T_10_1(),
      .F2Adef_T_10_2(),
      .F2Adef_T_10_3(),
      .F2Adef_T_10_4(),
      .F2Adef_T_10_5(),
      .F2Adef_T_10_6(),
      .F2Adef_T_11_0(),
      .F2Adef_T_11_1(),
      .F2Adef_T_11_2(),
      .F2Adef_T_11_3(),
      .F2Adef_T_12_0(),
      .F2Adef_T_12_1(),
      .F2Adef_T_12_2(),
      .F2Adef_T_12_3(),
      .F2Adef_T_12_4(),
      .F2Adef_T_12_5(),
      .F2Adef_T_12_6(),
      .F2Adef_T_13_0(),
      .F2Adef_T_13_1(),
      .F2Adef_T_13_2(),
      .F2Adef_T_13_3(),
      .F2Adef_T_14_0(),
      .F2Adef_T_14_1(),
      .F2Adef_T_14_2(),
      .F2Adef_T_14_3(),
      .F2Adef_T_14_4(),
      .F2Adef_T_14_5(),
      .F2Adef_T_14_6(),
      .F2Adef_T_15_0(),
      .F2Adef_T_15_1(),
      .F2Adef_T_15_2(),
      .F2Adef_T_15_3(),
      .F2Adef_T_16_0(),
      .F2Adef_T_16_1(),
      .F2Adef_T_16_2(),
      .F2Adef_T_16_3(),
      .F2Adef_T_16_4(),
      .F2Adef_T_16_5(),
      .F2Adef_T_16_6(),
      .F2Adef_T_17_0(tcdm_clk_p2_def),
      .F2Adef_T_17_1(),
      .F2Adef_T_17_2(),
      .F2Adef_T_17_3(),
      .F2Adef_T_18_0(),
      .F2Adef_T_18_1(),
      .F2Adef_T_18_2(),
      .F2Adef_T_18_3(),
      .F2Adef_T_18_4(),
      .F2Adef_T_18_5(),
      .F2Adef_T_18_6(),
      .F2Adef_T_19_0(),
      .F2Adef_T_19_1(),
      .F2Adef_T_19_2(),
      .F2Adef_T_19_3(),
      .F2Adef_T_1_0(),
      .F2Adef_T_1_1(),
      .F2Adef_T_1_2(),
      .F2Adef_T_1_3(),
      .F2Adef_T_20_0(),
      .F2Adef_T_20_1(),
      .F2Adef_T_20_2(),
      .F2Adef_T_20_3(),
      .F2Adef_T_20_4(),
      .F2Adef_T_20_5(),
      .F2Adef_T_20_6(),
      .F2Adef_T_21_0(),
      .F2Adef_T_21_1(),
      .F2Adef_T_21_2(),
      .F2Adef_T_21_3(),
      .F2Adef_T_22_0(),
      .F2Adef_T_22_1(),
      .F2Adef_T_22_2(),
      .F2Adef_T_22_3(),
      .F2Adef_T_22_4(),
      .F2Adef_T_22_5(),
      .F2Adef_T_22_6(),
      .F2Adef_T_23_0(tcdm_clk_p3_def),
      .F2Adef_T_23_1(),
      .F2Adef_T_23_2(),
      .F2Adef_T_23_3(),
      .F2Adef_T_24_0(),
      .F2Adef_T_24_1(),
      .F2Adef_T_24_2(),
      .F2Adef_T_24_3(),
      .F2Adef_T_24_4(),
      .F2Adef_T_24_5(),
      .F2Adef_T_24_6(),
      .F2Adef_T_25_0(),
      .F2Adef_T_25_1(),
      .F2Adef_T_25_2(),
      .F2Adef_T_25_3(),
      .F2Adef_T_26_0(),
      .F2Adef_T_26_1(),
      .F2Adef_T_26_2(),
      .F2Adef_T_26_3(),
      .F2Adef_T_26_4(),
      .F2Adef_T_26_5(),
      .F2Adef_T_26_6(),
      .F2Adef_T_27_0(),
      .F2Adef_T_27_1(),
      .F2Adef_T_27_2(),
      .F2Adef_T_27_3(),
      .F2Adef_T_28_0(),
      .F2Adef_T_28_1(),
      .F2Adef_T_28_2(),
      .F2Adef_T_28_3(),
      .F2Adef_T_28_4(),
      .F2Adef_T_28_5(),
      .F2Adef_T_28_6(),
      .F2Adef_T_29_0(),
      .F2Adef_T_29_1(),
      .F2Adef_T_29_2(),
      .F2Adef_T_29_3(),
      .F2Adef_T_2_0(),
      .F2Adef_T_2_1(),
      .F2Adef_T_2_2(),
      .F2Adef_T_2_3(),
      .F2Adef_T_2_4(),
      .F2Adef_T_2_5(),
      .F2Adef_T_2_6(),
      .F2Adef_T_30_0(),
      .F2Adef_T_30_1(),
      .F2Adef_T_30_2(),
      .F2Adef_T_30_3(),
      .F2Adef_T_30_4(),
      .F2Adef_T_30_5(),
      .F2Adef_T_30_6(),
      .F2Adef_T_31_0(),
      .F2Adef_T_31_1(),
      .F2Adef_T_31_2(),
      .F2Adef_T_31_3(),
      .F2Adef_T_32_0(),
      .F2Adef_T_32_1(),
      .F2Adef_T_32_2(),
      .F2Adef_T_32_3(),
      .F2Adef_T_32_4(),
      .F2Adef_T_32_5(),
      .F2Adef_T_32_6(),
      .F2Adef_T_3_0(tcdm_clk_p0_def),
      .F2Adef_T_3_1(),
      .F2Adef_T_3_2(),
      .F2Adef_T_3_3(),
      .F2Adef_T_4_0(),
      .F2Adef_T_4_1(),
      .F2Adef_T_4_2(),
      .F2Adef_T_4_3(),
      .F2Adef_T_4_4(),
      .F2Adef_T_4_5(),
      .F2Adef_T_4_6(),
      .F2Adef_T_5_0(),
      .F2Adef_T_5_1(),
      .F2Adef_T_5_2(),
      .F2Adef_T_5_3(),
      .F2Adef_T_6_0(),
      .F2Adef_T_6_1(),
      .F2Adef_T_6_2(),
      .F2Adef_T_6_3(),
      .F2Adef_T_6_4(),
      .F2Adef_T_6_5(),
      .F2Adef_T_6_6(),
      .F2Adef_T_7_0(),
      .F2Adef_T_7_1(),
      .F2Adef_T_7_2(),
      .F2Adef_T_7_3(),
      .F2Adef_T_8_0(),
      .F2Adef_T_8_1(),
      .F2Adef_T_8_2(),
      .F2Adef_T_8_3(),
      .F2Adef_T_8_4(),
      .F2Adef_T_8_5(),
      .F2Adef_T_8_6(),
      .F2Adef_T_9_0(tcdm_clk_p1_def),
      .F2Adef_T_9_1(),
      .F2Adef_T_9_2(),
      .F2Adef_T_9_3(),
      .F2Adef_R_10_0(),
      .F2Adef_R_10_1(),
      .F2Adef_R_10_2(),
      .F2Adef_R_10_3(),
      .F2Adef_R_10_4(),
      .F2Adef_R_10_5(),
      .F2Adef_R_10_6(),
      .F2Adef_R_11_0(),
      .F2Adef_R_11_1(),
      .F2Adef_R_11_2(),
      .F2Adef_R_11_3(),
      .F2Adef_R_12_0(),
      .F2Adef_R_12_1(),
      .F2Adef_R_12_2(),
      .F2Adef_R_12_3(),
      .F2Adef_R_12_4(),
      .F2Adef_R_12_5(),
      .F2Adef_R_12_6(),
      .F2Adef_R_13_0(m0_coef_powerdn),
      .F2Adef_R_13_1(m0_coef_wclk_def),
      .F2Adef_R_13_2(),
      .F2Adef_R_13_3(),
      .F2Adef_R_14_0(),
      .F2Adef_R_14_1(),
      .F2Adef_R_14_2(),
      .F2Adef_R_14_3(),
      .F2Adef_R_14_4(),
      .F2Adef_R_14_5(),
      .F2Adef_R_14_6(),
      .F2Adef_R_15_0(m0_coef_rclk_def),
      .F2Adef_R_15_1(),
      .F2Adef_R_15_2(),
      .F2Adef_R_15_3(),
      .F2Adef_R_16_0(),
      .F2Adef_R_16_1(),
      .F2Adef_R_16_2(),
      .F2Adef_R_16_3(),
      .F2Adef_R_16_4(),
      .F2Adef_R_16_5(),
      .F2Adef_R_16_6(),
      .F2Adef_R_17_0(),
      .F2Adef_R_17_1(),
      .F2Adef_R_17_2(),
      .F2Adef_R_17_3(),
      .F2Adef_R_18_0(),
      .F2Adef_R_18_1(),
      .F2Adef_R_18_2(),
      .F2Adef_R_18_3(),
      .F2Adef_R_18_4(),
      .F2Adef_R_18_5(),
      .F2Adef_R_18_6(),
      .F2Adef_R_19_0(m0_m1_clk_def),
      .F2Adef_R_19_1(),
      .F2Adef_R_19_2(),
      .F2Adef_R_19_3(),
      .F2Adef_R_1_0(),
      .F2Adef_R_1_1(),
      .F2Adef_R_1_2(),
      .F2Adef_R_1_3(),
      .F2Adef_R_20_0(),
      .F2Adef_R_20_1(),
      .F2Adef_R_20_2(),
      .F2Adef_R_20_3(),
      .F2Adef_R_20_4(),
      .F2Adef_R_20_5(),
      .F2Adef_R_20_6(),
      .F2Adef_R_21_0(),
      .F2Adef_R_21_1(),
      .F2Adef_R_21_2(),
      .F2Adef_R_21_3(),
      .F2Adef_R_22_0(),
      .F2Adef_R_22_1(),
      .F2Adef_R_22_2(),
      .F2Adef_R_22_3(),
      .F2Adef_R_22_4(),
      .F2Adef_R_22_5(),
      .F2Adef_R_22_6(),
      .F2Adef_R_23_0(),
      .F2Adef_R_23_1(),
      .F2Adef_R_23_2(),
      .F2Adef_R_23_3(),
      .F2Adef_R_24_0(m0_oper1_powerdn),
      .F2Adef_R_24_1(),
      .F2Adef_R_24_2(),
      .F2Adef_R_24_3(),
      .F2Adef_R_24_4(),
      .F2Adef_R_24_5(),
      .F2Adef_R_24_6(),
      .F2Adef_R_25_0(),
      .F2Adef_R_25_1(),
      .F2Adef_R_25_2(),
      .F2Adef_R_25_3(),
      .F2Adef_R_26_0(),
      .F2Adef_R_26_1(),
      .F2Adef_R_26_2(),
      .F2Adef_R_26_3(),
      .F2Adef_R_26_4(),
      .F2Adef_R_26_5(),
      .F2Adef_R_26_6(),
      .F2Adef_R_27_0(),
      .F2Adef_R_27_1(),
      .F2Adef_R_27_2(),
      .F2Adef_R_27_3(),
      .F2Adef_R_28_0(m0_oper1_wclk_def),
      .F2Adef_R_28_1(),
      .F2Adef_R_28_2(),
      .F2Adef_R_28_3(),
      .F2Adef_R_28_4(),
      .F2Adef_R_28_5(),
      .F2Adef_R_28_6(),
      .F2Adef_R_29_0(m0_oper1_rclk_def),
      .F2Adef_R_29_1(),
      .F2Adef_R_29_2(),
      .F2Adef_R_29_3(),
      .F2Adef_R_2_0(m0_oper0_wclk_def),
      .F2Adef_R_2_1(),
      .F2Adef_R_2_2(),
      .F2Adef_R_2_3(),
      .F2Adef_R_2_4(),
      .F2Adef_R_2_5(),
      .F2Adef_R_2_6(),
      .F2Adef_R_30_0(),
      .F2Adef_R_30_1(),
      .F2Adef_R_30_2(),
      .F2Adef_R_30_3(),
      .F2Adef_R_30_4(),
      .F2Adef_R_30_5(),
      .F2Adef_R_30_6(),
      .F2Adef_R_31_0(),
      .F2Adef_R_31_1(),
      .F2Adef_R_31_2(),
      .F2Adef_R_31_3(),
      .F2Adef_R_32_0(),
      .F2Adef_R_32_1(),
      .F2Adef_R_32_2(),
      .F2Adef_R_32_3(),
      .F2Adef_R_32_4(),
      .F2Adef_R_32_5(),
      .F2Adef_R_32_6(),
      .F2Adef_R_3_0(),
      .F2Adef_R_3_1(),
      .F2Adef_R_3_2(),
      .F2Adef_R_3_3(),
      .F2Adef_R_4_0(),
      .F2Adef_R_4_1(),
      .F2Adef_R_4_2(),
      .F2Adef_R_4_3(),
      .F2Adef_R_4_4(),
      .F2Adef_R_4_5(),
      .F2Adef_R_4_6(),
      .F2Adef_R_5_0(),
      .F2Adef_R_5_1(),
      .F2Adef_R_5_2(),
      .F2Adef_R_5_3(),
      .F2Adef_R_6_0(m0_oper0_rclk_def),
      .F2Adef_R_6_1(m0_oper0_powerdn),
      .F2Adef_R_6_2(),
      .F2Adef_R_6_3(),
      .F2Adef_R_6_4(),
      .F2Adef_R_6_5(),
      .F2Adef_R_6_6(),
      .F2Adef_R_7_0(m0_m0_clk_def),
      .F2Adef_R_7_1(),
      .F2Adef_R_7_2(),
      .F2Adef_R_7_3(),
      .F2Adef_R_8_0(),
      .F2Adef_R_8_1(),
      .F2Adef_R_8_2(),
      .F2Adef_R_8_3(),
      .F2Adef_R_8_4(),
      .F2Adef_R_8_5(),
      .F2Adef_R_8_6(),
      .F2Adef_R_9_0(),
      .F2Adef_R_9_1(),
      .F2Adef_R_9_2(),
      .F2Adef_R_9_3(),
      .F2Areg_B_11_0(),
      .F2Areg_B_11_1(),
      .F2Areg_B_13_0(),
      .F2Areg_B_13_1(),
      .F2Areg_B_15_0(),
      .F2Areg_B_15_1(),
      .F2Areg_B_17_0(),
      .F2Areg_B_17_1(),
      .F2Areg_B_19_0(),
      .F2Areg_B_19_1(),
      .F2Areg_B_1_0(),
      .F2Areg_B_1_1(),
      .F2Areg_B_21_0(),
      .F2Areg_B_21_1(),
      .F2Areg_B_23_0(),
      .F2Areg_B_23_1(),
      .F2Areg_B_25_0(),
      .F2Areg_B_25_1(),
      .F2Areg_B_27_0(),
      .F2Areg_B_27_1(),
      .F2Areg_B_29_0(),
      .F2Areg_B_29_1(),
      .F2Areg_B_31_0(),
      .F2Areg_B_31_1(),
      .F2Areg_B_3_0(),
      .F2Areg_B_3_1(),
      .F2Areg_B_5_0(),
      .F2Areg_B_5_1(),
      .F2Areg_B_7_0(),
      .F2Areg_B_7_1(),
      .F2Areg_B_9_0(),
      .F2Areg_B_9_1(),
      .F2Areg_L_11_0(),
      .F2Areg_L_11_1(),
      .F2Areg_L_13_0(),
      .F2Areg_L_13_1(),
      .F2Areg_L_15_0(),
      .F2Areg_L_15_1(),
      .F2Areg_L_17_0(),
      .F2Areg_L_17_1(),
      .F2Areg_L_19_0(),
      .F2Areg_L_19_1(),
      .F2Areg_L_1_0(),
      .F2Areg_L_1_1(),
      .F2Areg_L_21_0(),
      .F2Areg_L_21_1(),
      .F2Areg_L_23_0(),
      .F2Areg_L_23_1(),
      .F2Areg_L_25_0(),
      .F2Areg_L_25_1(),
      .F2Areg_L_27_0(),
      .F2Areg_L_27_1(),
      .F2Areg_L_29_0(),
      .F2Areg_L_29_1(),
      .F2Areg_L_31_0(),
      .F2Areg_L_31_1(),
      .F2Areg_L_3_0(),
      .F2Areg_L_3_1(),
      .F2Areg_L_5_0(),
      .F2Areg_L_5_1(),
      .F2Areg_L_7_0(),
      .F2Areg_L_7_1(),
      .F2Areg_L_9_0(),
      .F2Areg_L_9_1(),
      .F2Areg_T_11_0(),
      .F2Areg_T_11_1(),
      .F2Areg_T_13_0(),
      .F2Areg_T_13_1(),
      .F2Areg_T_15_0(),
      .F2Areg_T_15_1(),
      .F2Areg_T_17_0(),
      .F2Areg_T_17_1(),
      .F2Areg_T_19_0(),
      .F2Areg_T_19_1(),
      .F2Areg_T_1_0(),
      .F2Areg_T_1_1(),
      .F2Areg_T_21_0(),
      .F2Areg_T_21_1(),
      .F2Areg_T_23_0(),
      .F2Areg_T_23_1(),
      .F2Areg_T_25_0(),
      .F2Areg_T_25_1(),
      .F2Areg_T_27_0(),
      .F2Areg_T_27_1(),
      .F2Areg_T_29_0(),
      .F2Areg_T_29_1(),
      .F2Areg_T_31_0(),
      .F2Areg_T_31_1(),
      .F2Areg_T_3_0(),
      .F2Areg_T_3_1(),
      .F2Areg_T_5_0(),
      .F2Areg_T_5_1(),
      .F2Areg_T_7_0(),
      .F2Areg_T_7_1(),
      .F2Areg_T_9_0(),
      .F2Areg_T_9_1(),
      .F2Areg_R_11_0(),
      .F2Areg_R_11_1(),
      .F2Areg_R_13_0(),
      .F2Areg_R_13_1(),
      .F2Areg_R_15_0(),
      .F2Areg_R_15_1(),
      .F2Areg_R_17_0(),
      .F2Areg_R_17_1(),
      .F2Areg_R_19_0(),
      .F2Areg_R_19_1(),
      .F2Areg_R_1_0(),
      .F2Areg_R_1_1(),
      .F2Areg_R_21_0(),
      .F2Areg_R_21_1(),
      .F2Areg_R_23_0(),
      .F2Areg_R_23_1(),
      .F2Areg_R_25_0(),
      .F2Areg_R_25_1(),
      .F2Areg_R_27_0(),
      .F2Areg_R_27_1(),
      .F2Areg_R_29_0(),
      .F2Areg_R_29_1(),
      .F2Areg_R_31_0(),
      .F2Areg_R_31_1(),
      .F2Areg_R_3_0(),
      .F2Areg_R_3_1(),
      .F2Areg_R_5_0(),
      .F2Areg_R_5_1(),
      .F2Areg_R_7_0(),
      .F2Areg_R_7_1(),
      .F2Areg_R_9_0(),
      .F2Areg_R_9_1(),
      .BL_DOUT_0_(fcb_bl_dout[0]),
      .BL_DOUT_10_(fcb_bl_dout[10]),
      .BL_DOUT_11_(fcb_bl_dout[11]),
      .BL_DOUT_12_(fcb_bl_dout[12]),
      .BL_DOUT_13_(fcb_bl_dout[13]),
      .BL_DOUT_14_(fcb_bl_dout[14]),
      .BL_DOUT_15_(fcb_bl_dout[15]),
      .BL_DOUT_16_(fcb_bl_dout[16]),
      .BL_DOUT_17_(fcb_bl_dout[17]),
      .BL_DOUT_18_(fcb_bl_dout[18]),
      .BL_DOUT_19_(fcb_bl_dout[19]),
      .BL_DOUT_1_(fcb_bl_dout[1]),
      .BL_DOUT_20_(fcb_bl_dout[20]),
      .BL_DOUT_21_(fcb_bl_dout[21]),
      .BL_DOUT_22_(fcb_bl_dout[22]),
      .BL_DOUT_23_(fcb_bl_dout[23]),
      .BL_DOUT_24_(fcb_bl_dout[24]),
      .BL_DOUT_25_(fcb_bl_dout[25]),
      .BL_DOUT_26_(fcb_bl_dout[26]),
      .BL_DOUT_27_(fcb_bl_dout[27]),
      .BL_DOUT_28_(fcb_bl_dout[28]),
      .BL_DOUT_29_(fcb_bl_dout[29]),
      .BL_DOUT_2_(fcb_bl_dout[2]),
      .BL_DOUT_30_(fcb_bl_dout[30]),
      .BL_DOUT_31_(fcb_bl_dout[31]),
      .BL_DOUT_3_(fcb_bl_dout[3]),
      .BL_DOUT_4_(fcb_bl_dout[4]),
      .BL_DOUT_5_(fcb_bl_dout[5]),
      .BL_DOUT_6_(fcb_bl_dout[6]),
      .BL_DOUT_7_(fcb_bl_dout[7]),
      .BL_DOUT_8_(fcb_bl_dout[8]),
      .BL_DOUT_9_(fcb_bl_dout[9]),
      .FB_SPE_OUT_0_(FB_SPE_OUT[0]),
      .FB_SPE_OUT_1_(FB_SPE_OUT[1]),
      .FB_SPE_OUT_2_(FB_SPE_OUT[2]),
      .FB_SPE_OUT_3_(FB_SPE_OUT[3]),
      .PARALLEL_CFG(fcb_pif_en)
  );

endmodule



