module a2_bootrom #(
    parameter ADDR_WIDTH = 32,
    parameter DATA_WIDTH = 32
) (
    input  logic                  CLK,
    input  logic                  CEN,
    input  logic [ADDR_WIDTH-1:0] A,
    output logic [DATA_WIDTH-1:0] Q
);
  logic [31:0] value;
  assign Q = value;
  always @(posedge CLK) begin
    case (A)
      0: value <= 32'h09C0006F;
      1: value <= 32'h0980006F;
      2: value <= 32'h0940006F;
      3: value <= 32'h0900006F;
      4: value <= 32'h08C0006F;
      5: value <= 32'h0880006F;
      6: value <= 32'h0840006F;
      7: value <= 32'h0800006F;
      8: value <= 32'h07C0006F;
      9: value <= 32'h0780006F;
      10: value <= 32'h0740006F;
      11: value <= 32'h0700006F;
      12: value <= 32'h06C0006F;
      13: value <= 32'h0680006F;
      14: value <= 32'h0640006F;
      15: value <= 32'h0600006F;
      16: value <= 32'h05C0006F;
      17: value <= 32'h0580006F;
      18: value <= 32'h0540006F;
      19: value <= 32'h0500006F;
      20: value <= 32'h04C0006F;
      21: value <= 32'h0480006F;
      22: value <= 32'h0440006F;
      23: value <= 32'h0400006F;
      24: value <= 32'h03C0006F;
      25: value <= 32'h0380006F;
      26: value <= 32'h0340006F;
      27: value <= 32'h0300006F;
      28: value <= 32'h02C0006F;
      29: value <= 32'h0280006F;
      30: value <= 32'h0240006F;
      31: value <= 32'h0200006F;
      32: value <= 32'h0080006F;
      33: value <= 32'h0000006F;
      34: value <= 32'h0207E117;
      35: value <= 32'hCE410113;
      36: value <= 32'h1F00006F;
      37: value <= 32'h00060113;
      38: value <= 32'h00058067;
      39: value <= 32'h30200073;
      40: value <= 32'hCA09832A;
      41: value <= 32'h00058383;
      42: value <= 32'h00730023;
      43: value <= 32'h0305167D;
      44: value <= 32'hFA6D0585;
      45: value <= 32'h11018082;
      46: value <= 32'h0070C62A;
      47: value <= 32'h45054585;
      48: value <= 32'h2B85CE06;
      49: value <= 32'h610540F2;
      50: value <= 32'h11418082;
      51: value <= 32'hC6064535;
      52: value <= 32'h40B237DD;
      53: value <= 32'h01414529;
      54: value <= 32'h47A9BFF9;
      55: value <= 32'h00F51363;
      56: value <= 32'hBFD1B7ED;
      57: value <= 32'hC4221141;
      58: value <= 32'h842AC606;
      59: value <= 32'h00040503;
      60: value <= 32'h40B2E509;
      61: value <= 32'h01414422;
      62: value <= 32'h37C58082;
      63: value <= 32'hB7FD0405;
      64: value <= 32'h00455793;
      65: value <= 32'h8BBD1141;
      66: value <= 32'hC606C422;
      67: value <= 32'h0713842A;
      68: value <= 32'h85130390;
      69: value <= 32'h54630307;
      70: value <= 32'h851300A7;
      71: value <= 32'h3F750577;
      72: value <= 32'h0513883D;
      73: value <= 32'h07930304;
      74: value <= 32'hD4630390;
      75: value <= 32'h051300A7;
      76: value <= 32'h44220574;
      77: value <= 32'h014140B2;
      78: value <= 32'h1141B74D;
      79: value <= 32'h842AC422;
      80: value <= 32'hC6068121;
      81: value <= 32'h85223F75;
      82: value <= 32'h40B24422;
      83: value <= 32'hBF4D0141;
      84: value <= 32'hC4221141;
      85: value <= 32'h8141842A;
      86: value <= 32'h37C5C606;
      87: value <= 32'h44228522;
      88: value <= 32'h014140B2;
      89: value <= 32'h1141BFD9;
      90: value <= 32'h6485C226;
      91: value <= 32'h40848593;
      92: value <= 32'h4641C422;
      93: value <= 32'h95AA842A;
      94: value <= 32'hC6064501;
      95: value <= 32'h265D94A2;
      96: value <= 32'h40C4A603;
      97: value <= 32'hCE6347BD;
      98: value <= 32'hCE1100C7;
      99: value <= 32'h85936585;
      100: value <= 32'h95A24185;
      101: value <= 32'h40B24422;
      102: value <= 32'h06124492;
      103: value <= 32'h01414541;
      104: value <= 32'h4641A651;
      105: value <= 32'h40B2B7E5;
      106: value <= 32'h44924422;
      107: value <= 32'h80820141;
      108: value <= 32'hD64E7139;
      109: value <= 32'hDA266985;
      110: value <= 32'hD05AD84A;
      111: value <= 32'h8493892A;
      112: value <= 32'h6B094189;
      113: value <= 32'hC86AD256;
      114: value <= 32'hDC22DE06;
      115: value <= 32'hCE5ED452;
      116: value <= 32'hCA66CC62;
      117: value <= 32'h94CAC66E;
      118: value <= 32'h4A813779;
      119: value <= 32'h9B4A99CA;
      120: value <= 32'h01000D37;
      121: value <= 32'h40C9A783;
      122: value <= 32'h02FAE363;
      123: value <= 32'h1A000537;
      124: value <= 32'h67C50513;
      125: value <= 32'hA5033DC5;
      126: value <= 32'h3F994109;
      127: value <= 32'h1A000537;
      128: value <= 32'h67850513;
      129: value <= 32'hA78335C5;
      130: value <= 32'h97824109;
      131: value <= 32'h07B7A001;
      132: value <= 32'h85131A00;
      133: value <= 32'h35F96687;
      134: value <= 32'h3F1D8556;
      135: value <= 32'h1A0007B7;
      136: value <= 32'h68478513;
      137: value <= 32'h40C835C1;
      138: value <= 32'hE4000BB7;
      139: value <= 32'h370D4C01;
      140: value <= 32'h0044AA03;
      141: value <= 32'h0004AC83;
      142: value <= 32'h0084AD83;
      143: value <= 32'h44D49BD2;
      144: value <= 32'h00DC6563;
      145: value <= 32'h04C10A85;
      146: value <= 32'h2403BF71;
      147: value <= 32'hF563920B;
      148: value <= 32'h8413008D;
      149: value <= 32'h9871003D;
      150: value <= 32'hFB638622;
      151: value <= 32'h85D201AB;
      152: value <= 32'h24C98566;
      153: value <= 32'h9CA29A22;
      154: value <= 32'h408D8DB3;
      155: value <= 32'hBFC10C05;
      156: value <= 32'h856685CA;
      157: value <= 32'h86222C45;
      158: value <= 32'h855285CA;
      159: value <= 32'hB7DD3515;
      160: value <= 32'h1C0107B7;
      161: value <= 32'h65F1439C;
      162: value <= 32'h47B71101;
      163: value <= 32'h85931A10;
      164: value <= 32'h45052005;
      165: value <= 32'hCC22CE06;
      166: value <= 32'hA403CA26;
      167: value <= 32'hC84A0C47;
      168: value <= 32'h0537263D;
      169: value <= 32'h05131A00;
      170: value <= 32'h3D2D68C5;
      171: value <= 32'h85228805;
      172: value <= 32'h25B73545;
      173: value <= 32'h85930026;
      174: value <= 32'h45015A05;
      175: value <= 32'h458128F1;
      176: value <= 32'h2A694501;
      177: value <= 32'h45014581;
      178: value <= 32'h00282AE5;
      179: value <= 32'hE4092211;
      180: value <= 32'h02E00793;
      181: value <= 32'h00F10423;
      182: value <= 32'h000104A3;
      183: value <= 32'h4437EC19;
      184: value <= 32'h44851A10;
      185: value <= 32'h2A234905;
      186: value <= 32'h587C0724;
      187: value <= 32'h00978463;
      188: value <= 32'h3DB95868;
      189: value <= 32'h33FD0028;
      190: value <= 32'hC537B7FD;
      191: value <= 32'h67851C07;
      192: value <= 32'h00050413;
      193: value <= 32'h09336489;
      194: value <= 32'h05130094;
      195: value <= 32'h943E0005;
      196: value <= 32'h92F92023;
      197: value <= 32'h90092E23;
      198: value <= 32'h40042223;
      199: value <= 32'h92092223;
      200: value <= 32'h27833599;
      201: value <= 32'h28039209;
      202: value <= 32'hD73740C4;
      203: value <= 32'h88931C07;
      204: value <= 32'h06B3FFF7;
      205: value <= 32'h071340F0;
      206: value <= 32'h46014207;
      207: value <= 32'h1C000537;
      208: value <= 32'h92848493;
      209: value <= 32'h03061563;
      210: value <= 32'h97AA6789;
      211: value <= 32'hA0236605;
      212: value <= 32'h061392C7;
      213: value <= 32'h962A5196;
      214: value <= 32'h1A0005B7;
      215: value <= 32'h9007AE23;
      216: value <= 32'h9207A223;
      217: value <= 32'h40060613;
      218: value <= 32'h1B058593;
      219: value <= 32'h27833325;
      220: value <= 32'h6963FFC7;
      221: value <= 32'h430C00F5;
      222: value <= 32'h696395BE;
      223: value <= 32'h060500B5;
      224: value <= 32'hB7C90741;
      225: value <= 32'h009505B3;
      226: value <= 32'hFEB7FBE3;
      227: value <= 32'h97AE430C;
      228: value <= 32'hF53397C6;
      229: value <= 32'hB7E500D7;
      230: value <= 32'h1A102737;
      231: value <= 32'h47914714;
      232: value <= 32'h00A79533;
      233: value <= 32'hC7148EC9;
      234: value <= 32'h47934714;
      235: value <= 32'h8FF5FFF5;
      236: value <= 32'h431CC71C;
      237: value <= 32'h57B78D5D;
      238: value <= 32'h8793004C;
      239: value <= 32'hD7B3B407;
      240: value <= 32'hC30802B7;
      241: value <= 32'h1C07E737;
      242: value <= 32'h04234501;
      243: value <= 32'h808296F7;
      244: value <= 32'h1A102637;
      245: value <= 32'h18864703;
      246: value <= 32'h1C07E6B7;
      247: value <= 32'h18060793;
      248: value <= 32'h04239B3D;
      249: value <= 32'h470318E6;
      250: value <= 32'h9B3D1986;
      251: value <= 32'h18E60C23;
      252: value <= 32'h1A864703;
      253: value <= 32'h04239B3D;
      254: value <= 32'hC6831AE6;
      255: value <= 32'hE7379686;
      256: value <= 32'h07131C07;
      257: value <= 32'hC3149287;
      258: value <= 32'h100006B7;
      259: value <= 32'h06B7C354;
      260: value <= 32'h86932007;
      261: value <= 32'hC71409F6;
      262: value <= 32'h704706B7;
      263: value <= 32'hC754068D;
      264: value <= 32'h900006B7;
      265: value <= 32'hCB140685;
      266: value <= 32'h18A62023;
      267: value <= 32'hC3D44691;
      268: value <= 32'h18864683;
      269: value <= 32'h0106E693;
      270: value <= 32'h18D60423;
      271: value <= 32'h4751D398;
      272: value <= 32'h4703D3D8;
      273: value <= 32'h67131A86;
      274: value <= 32'h04230107;
      275: value <= 32'h27371AE6;
      276: value <= 32'h07931A10;
      277: value <= 32'h43DC1807;
      278: value <= 32'h8082FFED;
      279: value <= 32'h003427B7;
      280: value <= 32'h04378793;
      281: value <= 32'h051E953E;
      282: value <= 32'h02854783;
      283: value <= 32'h1C07E737;
      284: value <= 32'h96874703;
      285: value <= 32'h04239BBD;
      286: value <= 32'h478302F5;
      287: value <= 32'hE7930285;
      288: value <= 32'h04230207;
      289: value <= 32'hE7B702F5;
      290: value <= 32'h87931C07;
      291: value <= 32'hC3989287;
      292: value <= 32'h10000737;
      293: value <= 32'h07378DD9;
      294: value <= 32'h07132007;
      295: value <= 32'hC7980667;
      296: value <= 32'h90000737;
      297: value <= 32'hD11C0705;
      298: value <= 32'hC7D8C3CC;
      299: value <= 32'hD15C47C1;
      300: value <= 32'h02854783;
      301: value <= 32'h0107E793;
      302: value <= 32'h02F50423;
      303: value <= 32'h80824501;
      304: value <= 32'h003427B7;
      305: value <= 32'h04378793;
      306: value <= 32'h051E953E;
      307: value <= 32'h02854783;
      308: value <= 32'h1C07E737;
      309: value <= 32'h96874703;
      310: value <= 32'h04239BBD;
      311: value <= 32'h478302F5;
      312: value <= 32'hE7930285;
      313: value <= 32'h04230207;
      314: value <= 32'hE7B702F5;
      315: value <= 32'h87931C07;
      316: value <= 32'hC3989287;
      317: value <= 32'h10000737;
      318: value <= 32'h07378DD9;
      319: value <= 32'h07132007;
      320: value <= 32'hC7980997;
      321: value <= 32'h90000737;
      322: value <= 32'hD11C0705;
      323: value <= 32'hC7D8C3CC;
      324: value <= 32'hD15C47C1;
      325: value <= 32'h02854783;
      326: value <= 32'h0107E793;
      327: value <= 32'h02F50423;
      328: value <= 32'h80824501;
      329: value <= 32'h1A102837;
      330: value <= 32'h18884703;
      331: value <= 32'h1C07E6B7;
      332: value <= 32'h200708B7;
      333: value <= 32'h04239B3D;
      334: value <= 32'h470318E8;
      335: value <= 32'h03371988;
      336: value <= 32'h0793200F;
      337: value <= 32'h9B3D1808;
      338: value <= 32'h18E80C23;
      339: value <= 32'h1A884703;
      340: value <= 32'h04239B3D;
      341: value <= 32'hC6831AE8;
      342: value <= 32'hE7379686;
      343: value <= 32'h07131C07;
      344: value <= 32'hC3149287;
      345: value <= 32'h100006B7;
      346: value <= 32'h8693C354;
      347: value <= 32'hC7140038;
      348: value <= 32'h00855693;
      349: value <= 32'h82C106C2;
      350: value <= 32'h0FF57513;
      351: value <= 32'h0066E6B3;
      352: value <= 32'h01156533;
      353: value <= 32'hCB08C754;
      354: value <= 32'hFFF60693;
      355: value <= 32'h70470537;
      356: value <= 32'hCB548EC9;
      357: value <= 32'h900006B7;
      358: value <= 32'hCF140685;
      359: value <= 32'h18B82023;
      360: value <= 32'h4683C3D0;
      361: value <= 32'hE6931888;
      362: value <= 32'h04230106;
      363: value <= 32'hD39818D8;
      364: value <= 32'hD3D84771;
      365: value <= 32'h1A884703;
      366: value <= 32'h01076713;
      367: value <= 32'h1AE80423;
      368: value <= 32'h1A102737;
      369: value <= 32'h18070793;
      370: value <= 32'hFFED43DC;
      371: value <= 32'h27378082;
      372: value <= 32'h47141A10;
      373: value <= 32'h97B34785;
      374: value <= 32'h8EDD00A7;
      375: value <= 32'h4710C714;
      376: value <= 32'hFFF7C693;
      377: value <= 32'hC7148EF1;
      378: value <= 32'h8FD54314;
      379: value <= 32'h27B7C31C;
      380: value <= 32'h87930034;
      381: value <= 32'h953E0417;
      382: value <= 32'h004C57B7;
      383: value <= 32'hB4078793;
      384: value <= 32'h02B7D7B3;
      385: value <= 32'h07C2051E;
      386: value <= 32'h132383C1;
      387: value <= 32'h515C02F5;
      388: value <= 32'h0067E793;
      389: value <= 32'h515CD15C;
      390: value <= 32'h0107E793;
      391: value <= 32'h515CD15C;
      392: value <= 32'h1007E793;
      393: value <= 32'h515CD15C;
      394: value <= 32'h2007E793;
      395: value <= 32'h4501D15C;
      396: value <= 32'h27B78082;
      397: value <= 32'h87930034;
      398: value <= 32'h953E0417;
      399: value <= 32'h00751793;
      400: value <= 32'h4BD84501;
      401: value <= 32'hCB90EF11;
      402: value <= 32'hC703CBCC;
      403: value <= 32'h67130187;
      404: value <= 32'h8C230107;
      405: value <= 32'h4BD800E7;
      406: value <= 32'h0542E711;
      407: value <= 32'h80828141;
      408: value <= 32'hB7C50505;
      409: value <= 32'hBFC50505;
      410: value <= 32'h616F4C0A;
      411: value <= 32'h676E6964;
      412: value <= 32'h63655320;
      413: value <= 32'h6E6F6974;
      414: value <= 32'h00000020;
      415: value <= 32'h6D754A0A;
      416: value <= 32'h676E6970;
      417: value <= 32'h206F7420;
      418: value <= 32'h00000000;
      419: value <= 32'h2032410A;
      420: value <= 32'h746F6F42;
      421: value <= 32'h64616F6C;
      422: value <= 32'h42207265;
      423: value <= 32'h73746F6F;
      424: value <= 32'h003D6C65;
      425: value <= 32'h00000000;
      426: value <= 32'h00000000;
      427: value <= 32'h00000000;
      428: value <= 32'h00000000;
      429: value <= 32'h00000000;
      430: value <= 32'h00000000;
      431: value <= 32'h00000000;
      432: value <= 32'h00000000;
      433: value <= 32'h00000000;
      434: value <= 32'h00000000;
      435: value <= 32'h00000000;
      436: value <= 32'h00000000;
      437: value <= 32'h00000000;
      438: value <= 32'h00000000;
      439: value <= 32'h00000000;
      440: value <= 32'h00000000;
      441: value <= 32'h00000000;
      442: value <= 32'h00000000;
      443: value <= 32'h00000000;
      444: value <= 32'h00000000;
      445: value <= 32'h00000000;
      446: value <= 32'h00000000;
      447: value <= 32'h00000000;
      448: value <= 32'h00000000;
      449: value <= 32'h00000000;
      450: value <= 32'h00000000;
      451: value <= 32'h00000000;
      452: value <= 32'h00000000;
      453: value <= 32'h00000000;
      454: value <= 32'h00000000;
      455: value <= 32'h00000000;
      456: value <= 32'h00000000;
      457: value <= 32'h00000000;
      458: value <= 32'h00000000;
      459: value <= 32'h00000000;
      460: value <= 32'h00000000;
      461: value <= 32'h00000000;
      462: value <= 32'h00000000;
      463: value <= 32'h00000000;
      464: value <= 32'h00000000;
      465: value <= 32'h00000000;
      466: value <= 32'h00000000;
      467: value <= 32'h00000000;
      468: value <= 32'h00000000;
      469: value <= 32'h00000000;
      470: value <= 32'h00000000;
      471: value <= 32'h00000000;
      472: value <= 32'h00000000;
      473: value <= 32'h00000000;
      474: value <= 32'h00000000;
      475: value <= 32'h00000000;
      476: value <= 32'h00000000;
      477: value <= 32'h00000000;
      478: value <= 32'h00000000;
      479: value <= 32'h00000000;
      480: value <= 32'h00000000;
      481: value <= 32'h00000000;
      482: value <= 32'h00000000;
      483: value <= 32'h00000000;
      484: value <= 32'h00000000;
      485: value <= 32'h00000000;
      486: value <= 32'h00000000;
      487: value <= 32'h00000000;
      488: value <= 32'h00000000;
      489: value <= 32'h00000000;
      490: value <= 32'h00000000;
      491: value <= 32'h00000000;
      492: value <= 32'h00000000;
      493: value <= 32'h00000000;
      494: value <= 32'h00000000;
      495: value <= 32'h00000000;
      496: value <= 32'h00000000;
      497: value <= 32'h00000000;
      498: value <= 32'h00000000;
      499: value <= 32'h00000000;
      500: value <= 32'h00000000;
      501: value <= 32'h00000000;
      502: value <= 32'h00000000;
      503: value <= 32'h00000000;
      504: value <= 32'h00000000;
      505: value <= 32'h00000000;
      506: value <= 32'h00000000;
      507: value <= 32'h00000000;
      508: value <= 32'h00000000;
      509: value <= 32'h00000000;
      510: value <= 32'h00000000;
      511: value <= 32'h00000000;
      512: value <= 32'h00000000;
      513: value <= 32'h00000000;
      514: value <= 32'h00000000;
      515: value <= 32'h00000000;
      516: value <= 32'h00000000;
      517: value <= 32'h00000000;
      518: value <= 32'h00000000;
      519: value <= 32'h00000000;
      520: value <= 32'h00000000;
      521: value <= 32'h00000000;
      522: value <= 32'h00000000;
      523: value <= 32'h00000000;
      524: value <= 32'h00000000;
      525: value <= 32'h00000000;
      526: value <= 32'h00000000;
      527: value <= 32'h00000000;
      528: value <= 32'h00000000;
      529: value <= 32'h00000000;
      530: value <= 32'h00000000;
      531: value <= 32'h00000000;
      532: value <= 32'h00000000;
      533: value <= 32'h00000000;
      534: value <= 32'h00000000;
      535: value <= 32'h00000000;
      536: value <= 32'h00000000;
      537: value <= 32'h00000000;
      538: value <= 32'h00000000;
      539: value <= 32'h00000000;
      540: value <= 32'h00000000;
      541: value <= 32'h00000000;
      542: value <= 32'h00000000;
      543: value <= 32'h00000000;
      544: value <= 32'h00000000;
      545: value <= 32'h00000000;
      546: value <= 32'h00000000;
      547: value <= 32'h00000000;
      548: value <= 32'h00000000;
      549: value <= 32'h00000000;
      550: value <= 32'h00000000;
      551: value <= 32'h00000000;
      552: value <= 32'h00000000;
      553: value <= 32'h00000000;
      554: value <= 32'h00000000;
      555: value <= 32'h00000000;
      556: value <= 32'h00000000;
      557: value <= 32'h00000000;
      558: value <= 32'h00000000;
      559: value <= 32'h00000000;
      560: value <= 32'h00000000;
      561: value <= 32'h00000000;
      562: value <= 32'h00000000;
      563: value <= 32'h00000000;
      564: value <= 32'h00000000;
      565: value <= 32'h00000000;
      566: value <= 32'h00000000;
      567: value <= 32'h00000000;
      568: value <= 32'h00000000;
      569: value <= 32'h00000000;
      570: value <= 32'h00000000;
      571: value <= 32'h00000000;
      572: value <= 32'h00000000;
      573: value <= 32'h00000000;
      574: value <= 32'h00000000;
      575: value <= 32'h00000000;
      576: value <= 32'h00000000;
      577: value <= 32'h00000000;
      578: value <= 32'h00000000;
      579: value <= 32'h00000000;
      580: value <= 32'h00000000;
      581: value <= 32'h00000000;
      582: value <= 32'h00000000;
      583: value <= 32'h00000000;
      584: value <= 32'h00000000;
      585: value <= 32'h00000000;
      586: value <= 32'h00000000;
      587: value <= 32'h00000000;
      588: value <= 32'h00000000;
      589: value <= 32'h00000000;
      590: value <= 32'h00000000;
      591: value <= 32'h00000000;
      592: value <= 32'h00000000;
      593: value <= 32'h00000000;
      594: value <= 32'h00000000;
      595: value <= 32'h00000000;
      596: value <= 32'h00000000;
      597: value <= 32'h00000000;
      598: value <= 32'h00000000;
      599: value <= 32'h00000000;
      600: value <= 32'h00000000;
      601: value <= 32'h00000000;
      602: value <= 32'h00000000;
      603: value <= 32'h00000000;
      604: value <= 32'h00000000;
      605: value <= 32'h00000000;
      606: value <= 32'h00000000;
      607: value <= 32'h00000000;
      608: value <= 32'h00000000;
      609: value <= 32'h00000000;
      610: value <= 32'h00000000;
      611: value <= 32'h00000000;
      612: value <= 32'h00000000;
      613: value <= 32'h00000000;
      614: value <= 32'h00000000;
      615: value <= 32'h00000000;
      616: value <= 32'h00000000;
      617: value <= 32'h00000000;
      618: value <= 32'h00000000;
      619: value <= 32'h00000000;
      620: value <= 32'h00000000;
      621: value <= 32'h00000000;
      622: value <= 32'h00000000;
      623: value <= 32'h00000000;
      624: value <= 32'h00000000;
      625: value <= 32'h00000000;
      626: value <= 32'h00000000;
      627: value <= 32'h00000000;
      628: value <= 32'h00000000;
      629: value <= 32'h00000000;
      630: value <= 32'h00000000;
      631: value <= 32'h00000000;
      632: value <= 32'h00000000;
      633: value <= 32'h00000000;
      634: value <= 32'h00000000;
      635: value <= 32'h00000000;
      636: value <= 32'h00000000;
      637: value <= 32'h00000000;
      638: value <= 32'h00000000;
      639: value <= 32'h00000000;
      640: value <= 32'h00000000;
      641: value <= 32'h00000000;
      642: value <= 32'h00000000;
      643: value <= 32'h00000000;
      644: value <= 32'h00000000;
      645: value <= 32'h00000000;
      646: value <= 32'h00000000;
      647: value <= 32'h00000000;
      648: value <= 32'h00000000;
      649: value <= 32'h00000000;
      650: value <= 32'h00000000;
      651: value <= 32'h00000000;
      652: value <= 32'h00000000;
      653: value <= 32'h00000000;
      654: value <= 32'h00000000;
      655: value <= 32'h00000000;
      656: value <= 32'h00000000;
      657: value <= 32'h00000000;
      658: value <= 32'h00000000;
      659: value <= 32'h00000000;
      660: value <= 32'h00000000;
      661: value <= 32'h00000000;
      662: value <= 32'h00000000;
      663: value <= 32'h00000000;
      664: value <= 32'h00000000;
      665: value <= 32'h00000000;
      666: value <= 32'h00000000;
      667: value <= 32'h00000000;
      668: value <= 32'h00000000;
      669: value <= 32'h00000000;
      670: value <= 32'h00000000;
      671: value <= 32'h00000000;
      672: value <= 32'h00000000;
      673: value <= 32'h00000000;
      674: value <= 32'h00000000;
      675: value <= 32'h00000000;
      676: value <= 32'h00000000;
      677: value <= 32'h00000000;
      678: value <= 32'h00000000;
      679: value <= 32'h00000000;
      680: value <= 32'h00000000;
      681: value <= 32'h00000000;
      682: value <= 32'h00000000;
      683: value <= 32'h00000000;
      684: value <= 32'h00000000;
      685: value <= 32'h00000000;
      686: value <= 32'h00000000;
      687: value <= 32'h00000000;
      688: value <= 32'h00000000;
      689: value <= 32'h00000000;
      690: value <= 32'h00000000;
      691: value <= 32'h00000000;
      692: value <= 32'h00000000;
      693: value <= 32'h00000000;
      694: value <= 32'h00000000;
      695: value <= 32'h00000000;
      696: value <= 32'h00000000;
      697: value <= 32'h00000000;
      698: value <= 32'h00000000;
      699: value <= 32'h00000000;
      700: value <= 32'h00000000;
      701: value <= 32'h00000000;
      702: value <= 32'h00000000;
      703: value <= 32'h00000000;
      704: value <= 32'h00000000;
      705: value <= 32'h00000000;
      706: value <= 32'h00000000;
      707: value <= 32'h00000000;
      708: value <= 32'h00000000;
      709: value <= 32'h00000000;
      710: value <= 32'h00000000;
      711: value <= 32'h00000000;
      712: value <= 32'h00000000;
      713: value <= 32'h00000000;
      714: value <= 32'h00000000;
      715: value <= 32'h00000000;
      716: value <= 32'h00000000;
      717: value <= 32'h00000000;
      718: value <= 32'h00000000;
      719: value <= 32'h00000000;
      720: value <= 32'h00000000;
      721: value <= 32'h00000000;
      722: value <= 32'h00000000;
      723: value <= 32'h00000000;
      724: value <= 32'h00000000;
      725: value <= 32'h00000000;
      726: value <= 32'h00000000;
      727: value <= 32'h00000000;
      728: value <= 32'h00000000;
      729: value <= 32'h00000000;
      730: value <= 32'h00000000;
      731: value <= 32'h00000000;
      732: value <= 32'h00000000;
      733: value <= 32'h00000000;
      734: value <= 32'h00000000;
      735: value <= 32'h00000000;
      736: value <= 32'h00000000;
      737: value <= 32'h00000000;
      738: value <= 32'h00000000;
      739: value <= 32'h00000000;
      740: value <= 32'h00000000;
      741: value <= 32'h00000000;
      742: value <= 32'h00000000;
      743: value <= 32'h00000000;
      744: value <= 32'h00000000;
      745: value <= 32'h00000000;
      746: value <= 32'h00000000;
      747: value <= 32'h00000000;
      748: value <= 32'h00000000;
      749: value <= 32'h00000000;
      750: value <= 32'h00000000;
      751: value <= 32'h00000000;
      752: value <= 32'h00000000;
      753: value <= 32'h00000000;
      754: value <= 32'h00000000;
      755: value <= 32'h00000000;
      756: value <= 32'h00000000;
      757: value <= 32'h00000000;
      758: value <= 32'h00000000;
      759: value <= 32'h00000000;
      760: value <= 32'h00000000;
      761: value <= 32'h00000000;
      762: value <= 32'h00000000;
      763: value <= 32'h00000000;
      764: value <= 32'h00000000;
      765: value <= 32'h00000000;
      766: value <= 32'h00000000;
      767: value <= 32'h00000000;
      768: value <= 32'h00000000;
      769: value <= 32'h00000000;
      770: value <= 32'h00000000;
      771: value <= 32'h00000000;
      772: value <= 32'h00000000;
      773: value <= 32'h00000000;
      774: value <= 32'h00000000;
      775: value <= 32'h00000000;
      776: value <= 32'h00000000;
      777: value <= 32'h00000000;
      778: value <= 32'h00000000;
      779: value <= 32'h00000000;
      780: value <= 32'h00000000;
      781: value <= 32'h00000000;
      782: value <= 32'h00000000;
      783: value <= 32'h00000000;
      784: value <= 32'h00000000;
      785: value <= 32'h00000000;
      786: value <= 32'h00000000;
      787: value <= 32'h00000000;
      788: value <= 32'h00000000;
      789: value <= 32'h00000000;
      790: value <= 32'h00000000;
      791: value <= 32'h00000000;
      792: value <= 32'h00000000;
      793: value <= 32'h00000000;
      794: value <= 32'h00000000;
      795: value <= 32'h00000000;
      796: value <= 32'h00000000;
      797: value <= 32'h00000000;
      798: value <= 32'h00000000;
      799: value <= 32'h00000000;
      800: value <= 32'h00000000;
      801: value <= 32'h00000000;
      802: value <= 32'h00000000;
      803: value <= 32'h00000000;
      804: value <= 32'h00000000;
      805: value <= 32'h00000000;
      806: value <= 32'h00000000;
      807: value <= 32'h00000000;
      808: value <= 32'h00000000;
      809: value <= 32'h00000000;
      810: value <= 32'h00000000;
      811: value <= 32'h00000000;
      812: value <= 32'h00000000;
      813: value <= 32'h00000000;
      814: value <= 32'h00000000;
      815: value <= 32'h00000000;
      816: value <= 32'h00000000;
      817: value <= 32'h00000000;
      818: value <= 32'h00000000;
      819: value <= 32'h00000000;
      820: value <= 32'h00000000;
      821: value <= 32'h00000000;
      822: value <= 32'h00000000;
      823: value <= 32'h00000000;
      824: value <= 32'h00000000;
      825: value <= 32'h00000000;
      826: value <= 32'h00000000;
      827: value <= 32'h00000000;
      828: value <= 32'h00000000;
      829: value <= 32'h00000000;
      830: value <= 32'h00000000;
      831: value <= 32'h00000000;
      832: value <= 32'h00000000;
      833: value <= 32'h00000000;
      834: value <= 32'h00000000;
      835: value <= 32'h00000000;
      836: value <= 32'h00000000;
      837: value <= 32'h00000000;
      838: value <= 32'h00000000;
      839: value <= 32'h00000000;
      840: value <= 32'h00000000;
      841: value <= 32'h00000000;
      842: value <= 32'h00000000;
      843: value <= 32'h00000000;
      844: value <= 32'h00000000;
      845: value <= 32'h00000000;
      846: value <= 32'h00000000;
      847: value <= 32'h00000000;
      848: value <= 32'h00000000;
      849: value <= 32'h00000000;
      850: value <= 32'h00000000;
      851: value <= 32'h00000000;
      852: value <= 32'h00000000;
      853: value <= 32'h00000000;
      854: value <= 32'h00000000;
      855: value <= 32'h00000000;
      856: value <= 32'h00000000;
      857: value <= 32'h00000000;
      858: value <= 32'h00000000;
      859: value <= 32'h00000000;
      860: value <= 32'h00000000;
      861: value <= 32'h00000000;
      862: value <= 32'h00000000;
      863: value <= 32'h00000000;
      864: value <= 32'h00000000;
      865: value <= 32'h00000000;
      866: value <= 32'h00000000;
      867: value <= 32'h00000000;
      868: value <= 32'h00000000;
      869: value <= 32'h00000000;
      870: value <= 32'h00000000;
      871: value <= 32'h00000000;
      872: value <= 32'h00000000;
      873: value <= 32'h00000000;
      874: value <= 32'h00000000;
      875: value <= 32'h00000000;
      876: value <= 32'h00000000;
      877: value <= 32'h00000000;
      878: value <= 32'h00000000;
      879: value <= 32'h00000000;
      880: value <= 32'h00000000;
      881: value <= 32'h00000000;
      882: value <= 32'h00000000;
      883: value <= 32'h00000000;
      884: value <= 32'h00000000;
      885: value <= 32'h00000000;
      886: value <= 32'h00000000;
      887: value <= 32'h00000000;
      888: value <= 32'h00000000;
      889: value <= 32'h00000000;
      890: value <= 32'h00000000;
      891: value <= 32'h00000000;
      892: value <= 32'h00000000;
      893: value <= 32'h00000000;
      894: value <= 32'h00000000;
      895: value <= 32'h00000000;
      896: value <= 32'h00000000;
      897: value <= 32'h00000000;
      898: value <= 32'h00000000;
      899: value <= 32'h00000000;
      900: value <= 32'h00000000;
      901: value <= 32'h00000000;
      902: value <= 32'h00000000;
      903: value <= 32'h00000000;
      904: value <= 32'h00000000;
      905: value <= 32'h00000000;
      906: value <= 32'h00000000;
      907: value <= 32'h00000000;
      908: value <= 32'h00000000;
      909: value <= 32'h00000000;
      910: value <= 32'h00000000;
      911: value <= 32'h00000000;
      912: value <= 32'h00000000;
      913: value <= 32'h00000000;
      914: value <= 32'h00000000;
      915: value <= 32'h00000000;
      916: value <= 32'h00000000;
      917: value <= 32'h00000000;
      918: value <= 32'h00000000;
      919: value <= 32'h00000000;
      920: value <= 32'h00000000;
      921: value <= 32'h00000000;
      922: value <= 32'h00000000;
      923: value <= 32'h00000000;
      924: value <= 32'h00000000;
      925: value <= 32'h00000000;
      926: value <= 32'h00000000;
      927: value <= 32'h00000000;
      928: value <= 32'h00000000;
      929: value <= 32'h00000000;
      930: value <= 32'h00000000;
      931: value <= 32'h00000000;
      932: value <= 32'h00000000;
      933: value <= 32'h00000000;
      934: value <= 32'h00000000;
      935: value <= 32'h00000000;
      936: value <= 32'h00000000;
      937: value <= 32'h00000000;
      938: value <= 32'h00000000;
      939: value <= 32'h00000000;
      940: value <= 32'h00000000;
      941: value <= 32'h00000000;
      942: value <= 32'h00000000;
      943: value <= 32'h00000000;
      944: value <= 32'h00000000;
      945: value <= 32'h00000000;
      946: value <= 32'h00000000;
      947: value <= 32'h00000000;
      948: value <= 32'h00000000;
      949: value <= 32'h00000000;
      950: value <= 32'h00000000;
      951: value <= 32'h00000000;
      952: value <= 32'h00000000;
      953: value <= 32'h00000000;
      954: value <= 32'h00000000;
      955: value <= 32'h00000000;
      956: value <= 32'h00000000;
      957: value <= 32'h00000000;
      958: value <= 32'h00000000;
      959: value <= 32'h00000000;
      960: value <= 32'h00000000;
      961: value <= 32'h00000000;
      962: value <= 32'h00000000;
      963: value <= 32'h00000000;
      964: value <= 32'h00000000;
      965: value <= 32'h00000000;
      966: value <= 32'h00000000;
      967: value <= 32'h00000000;
      968: value <= 32'h00000000;
      969: value <= 32'h00000000;
      970: value <= 32'h00000000;
      971: value <= 32'h00000000;
      972: value <= 32'h00000000;
      973: value <= 32'h00000000;
      974: value <= 32'h00000000;
      975: value <= 32'h00000000;
      976: value <= 32'h00000000;
      977: value <= 32'h00000000;
      978: value <= 32'h00000000;
      979: value <= 32'h00000000;
      980: value <= 32'h00000000;
      981: value <= 32'h00000000;
      982: value <= 32'h00000000;
      983: value <= 32'h00000000;
      984: value <= 32'h00000000;
      985: value <= 32'h00000000;
      986: value <= 32'h00000000;
      987: value <= 32'h00000000;
      988: value <= 32'h00000000;
      989: value <= 32'h00000000;
      990: value <= 32'h00000000;
      991: value <= 32'h00000000;
      992: value <= 32'h00000000;
      993: value <= 32'h00000000;
      994: value <= 32'h00000000;
      995: value <= 32'h00000000;
      996: value <= 32'h00000000;
      997: value <= 32'h00000000;
      998: value <= 32'h00000000;
      999: value <= 32'h00000000;
      1000: value <= 32'h00000000;
      1001: value <= 32'h00000000;
      1002: value <= 32'h00000000;
      1003: value <= 32'h00000000;
      1004: value <= 32'h00000000;
      1005: value <= 32'h00000000;
      1006: value <= 32'h00000000;
      1007: value <= 32'h00000000;
      1008: value <= 32'h00000000;
      1009: value <= 32'h00000000;
      1010: value <= 32'h00000000;
      1011: value <= 32'h00000000;
      1012: value <= 32'h00000000;
      1013: value <= 32'h00000000;
      1014: value <= 32'h00000000;
      1015: value <= 32'h00000000;
      1016: value <= 32'h00000000;
      1017: value <= 32'h00000000;
      1018: value <= 32'h00000000;
      1019: value <= 32'h00000000;
      1020: value <= 32'h00000000;
      1021: value <= 32'h00000000;
      1022: value <= 32'h00000000;
      1023: value <= 32'h00000000;
      1024: value <= 32'h00000000;
      1025: value <= 32'h00000000;
      1026: value <= 32'h00000000;
      1027: value <= 32'h00000000;
      1028: value <= 32'h00000000;
      1029: value <= 32'h00000000;
      1030: value <= 32'h00000000;
      1031: value <= 32'h00000000;
      1032: value <= 32'h00000000;
      1033: value <= 32'h00000000;
      1034: value <= 32'h00000000;
      1035: value <= 32'h00000000;
      1036: value <= 32'h00000000;
      1037: value <= 32'h00000000;
      1038: value <= 32'h00000000;
      1039: value <= 32'h00000000;
      1040: value <= 32'h00000000;
      1041: value <= 32'h00000000;
      1042: value <= 32'h00000000;
      1043: value <= 32'h00000000;
      1044: value <= 32'h00000000;
      1045: value <= 32'h00000000;
      1046: value <= 32'h00000000;
      1047: value <= 32'h00000000;
      1048: value <= 32'h00000000;
      1049: value <= 32'h00000000;
      1050: value <= 32'h00000000;
      1051: value <= 32'h00000000;
      1052: value <= 32'h00000000;
      1053: value <= 32'h00000000;
      1054: value <= 32'h00000000;
      1055: value <= 32'h00000000;
      1056: value <= 32'h00000000;
      1057: value <= 32'h00000000;
      1058: value <= 32'h00000000;
      1059: value <= 32'h00000000;
      1060: value <= 32'h00000000;
      1061: value <= 32'h00000000;
      1062: value <= 32'h00000000;
      1063: value <= 32'h00000000;
      1064: value <= 32'h00000000;
      1065: value <= 32'h00000000;
      1066: value <= 32'h00000000;
      1067: value <= 32'h00000000;
      1068: value <= 32'h00000000;
      1069: value <= 32'h00000000;
      1070: value <= 32'h00000000;
      1071: value <= 32'h00000000;
      1072: value <= 32'h00000000;
      1073: value <= 32'h00000000;
      1074: value <= 32'h00000000;
      1075: value <= 32'h00000000;
      1076: value <= 32'h00000000;
      1077: value <= 32'h00000000;
      1078: value <= 32'h00000000;
      1079: value <= 32'h00000000;
      1080: value <= 32'h00000000;
      1081: value <= 32'h00000000;
      1082: value <= 32'h00000000;
      1083: value <= 32'h00000000;
      1084: value <= 32'h00000000;
      1085: value <= 32'h00000000;
      1086: value <= 32'h00000000;
      1087: value <= 32'h00000000;
      1088: value <= 32'h00000000;
      1089: value <= 32'h00000000;
      1090: value <= 32'h00000000;
      1091: value <= 32'h00000000;
      1092: value <= 32'h00000000;
      1093: value <= 32'h00000000;
      1094: value <= 32'h00000000;
      1095: value <= 32'h00000000;
      1096: value <= 32'h00000000;
      1097: value <= 32'h00000000;
      1098: value <= 32'h00000000;
      1099: value <= 32'h00000000;
      1100: value <= 32'h00000000;
      1101: value <= 32'h00000000;
      1102: value <= 32'h00000000;
      1103: value <= 32'h00000000;
      1104: value <= 32'h00000000;
      1105: value <= 32'h00000000;
      1106: value <= 32'h00000000;
      1107: value <= 32'h00000000;
      1108: value <= 32'h00000000;
      1109: value <= 32'h00000000;
      1110: value <= 32'h00000000;
      1111: value <= 32'h00000000;
      1112: value <= 32'h00000000;
      1113: value <= 32'h00000000;
      1114: value <= 32'h00000000;
      1115: value <= 32'h00000000;
      1116: value <= 32'h00000000;
      1117: value <= 32'h00000000;
      1118: value <= 32'h00000000;
      1119: value <= 32'h00000000;
      1120: value <= 32'h00000000;
      1121: value <= 32'h00000000;
      1122: value <= 32'h00000000;
      1123: value <= 32'h00000000;
      1124: value <= 32'h00000000;
      1125: value <= 32'h00000000;
      1126: value <= 32'h00000000;
      1127: value <= 32'h00000000;
      1128: value <= 32'h00000000;
      1129: value <= 32'h00000000;
      1130: value <= 32'h00000000;
      1131: value <= 32'h00000000;
      1132: value <= 32'h00000000;
      1133: value <= 32'h00000000;
      1134: value <= 32'h00000000;
      1135: value <= 32'h00000000;
      1136: value <= 32'h00000000;
      1137: value <= 32'h00000000;
      1138: value <= 32'h00000000;
      1139: value <= 32'h00000000;
      1140: value <= 32'h00000000;
      1141: value <= 32'h00000000;
      1142: value <= 32'h00000000;
      1143: value <= 32'h00000000;
      1144: value <= 32'h00000000;
      1145: value <= 32'h00000000;
      1146: value <= 32'h00000000;
      1147: value <= 32'h00000000;
      1148: value <= 32'h00000000;
      1149: value <= 32'h00000000;
      1150: value <= 32'h00000000;
      1151: value <= 32'h00000000;
      1152: value <= 32'h00000000;
      1153: value <= 32'h00000000;
      1154: value <= 32'h00000000;
      1155: value <= 32'h00000000;
      1156: value <= 32'h00000000;
      1157: value <= 32'h00000000;
      1158: value <= 32'h00000000;
      1159: value <= 32'h00000000;
      1160: value <= 32'h00000000;
      1161: value <= 32'h00000000;
      1162: value <= 32'h00000000;
      1163: value <= 32'h00000000;
      1164: value <= 32'h00000000;
      1165: value <= 32'h00000000;
      1166: value <= 32'h00000000;
      1167: value <= 32'h00000000;
      1168: value <= 32'h00000000;
      1169: value <= 32'h00000000;
      1170: value <= 32'h00000000;
      1171: value <= 32'h00000000;
      1172: value <= 32'h00000000;
      1173: value <= 32'h00000000;
      1174: value <= 32'h00000000;
      1175: value <= 32'h00000000;
      1176: value <= 32'h00000000;
      1177: value <= 32'h00000000;
      1178: value <= 32'h00000000;
      1179: value <= 32'h00000000;
      1180: value <= 32'h00000000;
      1181: value <= 32'h00000000;
      1182: value <= 32'h00000000;
      1183: value <= 32'h00000000;
      1184: value <= 32'h00000000;
      1185: value <= 32'h00000000;
      1186: value <= 32'h00000000;
      1187: value <= 32'h00000000;
      1188: value <= 32'h00000000;
      1189: value <= 32'h00000000;
      1190: value <= 32'h00000000;
      1191: value <= 32'h00000000;
      1192: value <= 32'h00000000;
      1193: value <= 32'h00000000;
      1194: value <= 32'h00000000;
      1195: value <= 32'h00000000;
      1196: value <= 32'h00000000;
      1197: value <= 32'h00000000;
      1198: value <= 32'h00000000;
      1199: value <= 32'h00000000;
      1200: value <= 32'h00000000;
      1201: value <= 32'h00000000;
      1202: value <= 32'h00000000;
      1203: value <= 32'h00000000;
      1204: value <= 32'h00000000;
      1205: value <= 32'h00000000;
      1206: value <= 32'h00000000;
      1207: value <= 32'h00000000;
      1208: value <= 32'h00000000;
      1209: value <= 32'h00000000;
      1210: value <= 32'h00000000;
      1211: value <= 32'h00000000;
      1212: value <= 32'h00000000;
      1213: value <= 32'h00000000;
      1214: value <= 32'h00000000;
      1215: value <= 32'h00000000;
      1216: value <= 32'h00000000;
      1217: value <= 32'h00000000;
      1218: value <= 32'h00000000;
      1219: value <= 32'h00000000;
      1220: value <= 32'h00000000;
      1221: value <= 32'h00000000;
      1222: value <= 32'h00000000;
      1223: value <= 32'h00000000;
      1224: value <= 32'h00000000;
      1225: value <= 32'h00000000;
      1226: value <= 32'h00000000;
      1227: value <= 32'h00000000;
      1228: value <= 32'h00000000;
      1229: value <= 32'h00000000;
      1230: value <= 32'h00000000;
      1231: value <= 32'h00000000;
      1232: value <= 32'h00000000;
      1233: value <= 32'h00000000;
      1234: value <= 32'h00000000;
      1235: value <= 32'h00000000;
      1236: value <= 32'h00000000;
      1237: value <= 32'h00000000;
      1238: value <= 32'h00000000;
      1239: value <= 32'h00000000;
      1240: value <= 32'h00000000;
      1241: value <= 32'h00000000;
      1242: value <= 32'h00000000;
      1243: value <= 32'h00000000;
      1244: value <= 32'h00000000;
      1245: value <= 32'h00000000;
      1246: value <= 32'h00000000;
      1247: value <= 32'h00000000;
      1248: value <= 32'h00000000;
      1249: value <= 32'h00000000;
      1250: value <= 32'h00000000;
      1251: value <= 32'h00000000;
      1252: value <= 32'h00000000;
      1253: value <= 32'h00000000;
      1254: value <= 32'h00000000;
      1255: value <= 32'h00000000;
      1256: value <= 32'h00000000;
      1257: value <= 32'h00000000;
      1258: value <= 32'h00000000;
      1259: value <= 32'h00000000;
      1260: value <= 32'h00000000;
      1261: value <= 32'h00000000;
      1262: value <= 32'h00000000;
      1263: value <= 32'h00000000;
      1264: value <= 32'h00000000;
      1265: value <= 32'h00000000;
      1266: value <= 32'h00000000;
      1267: value <= 32'h00000000;
      1268: value <= 32'h00000000;
      1269: value <= 32'h00000000;
      1270: value <= 32'h00000000;
      1271: value <= 32'h00000000;
      1272: value <= 32'h00000000;
      1273: value <= 32'h00000000;
      1274: value <= 32'h00000000;
      1275: value <= 32'h00000000;
      1276: value <= 32'h00000000;
      1277: value <= 32'h00000000;
      1278: value <= 32'h00000000;
      1279: value <= 32'h00000000;
      1280: value <= 32'h00000000;
      1281: value <= 32'h00000000;
      1282: value <= 32'h00000000;
      1283: value <= 32'h00000000;
      1284: value <= 32'h00000000;
      1285: value <= 32'h00000000;
      1286: value <= 32'h00000000;
      1287: value <= 32'h00000000;
      1288: value <= 32'h00000000;
      1289: value <= 32'h00000000;
      1290: value <= 32'h00000000;
      1291: value <= 32'h00000000;
      1292: value <= 32'h00000000;
      1293: value <= 32'h00000000;
      1294: value <= 32'h00000000;
      1295: value <= 32'h00000000;
      1296: value <= 32'h00000000;
      1297: value <= 32'h00000000;
      1298: value <= 32'h00000000;
      1299: value <= 32'h00000000;
      1300: value <= 32'h00000000;
      1301: value <= 32'h00000000;
      1302: value <= 32'h00000000;
      1303: value <= 32'h00000000;
      1304: value <= 32'h00000000;
      1305: value <= 32'h00000000;
      1306: value <= 32'h00000000;
      1307: value <= 32'h00000000;
      1308: value <= 32'h00000000;
      1309: value <= 32'h00000000;
      1310: value <= 32'h00000000;
      1311: value <= 32'h00000000;
      1312: value <= 32'h00000000;
      1313: value <= 32'h00000000;
      1314: value <= 32'h00000000;
      1315: value <= 32'h00000000;
      1316: value <= 32'h00000000;
      1317: value <= 32'h00000000;
      1318: value <= 32'h00000000;
      1319: value <= 32'h00000000;
      1320: value <= 32'h00000000;
      1321: value <= 32'h00000000;
      1322: value <= 32'h00000000;
      1323: value <= 32'h00000000;
      1324: value <= 32'h00000000;
      1325: value <= 32'h00000000;
      1326: value <= 32'h00000000;
      1327: value <= 32'h00000000;
      1328: value <= 32'h00000000;
      1329: value <= 32'h00000000;
      1330: value <= 32'h00000000;
      1331: value <= 32'h00000000;
      1332: value <= 32'h00000000;
      1333: value <= 32'h00000000;
      1334: value <= 32'h00000000;
      1335: value <= 32'h00000000;
      1336: value <= 32'h00000000;
      1337: value <= 32'h00000000;
      1338: value <= 32'h00000000;
      1339: value <= 32'h00000000;
      1340: value <= 32'h00000000;
      1341: value <= 32'h00000000;
      1342: value <= 32'h00000000;
      1343: value <= 32'h00000000;
      1344: value <= 32'h00000000;
      1345: value <= 32'h00000000;
      1346: value <= 32'h00000000;
      1347: value <= 32'h00000000;
      1348: value <= 32'h00000000;
      1349: value <= 32'h00000000;
      1350: value <= 32'h00000000;
      1351: value <= 32'h00000000;
      1352: value <= 32'h00000000;
      1353: value <= 32'h00000000;
      1354: value <= 32'h00000000;
      1355: value <= 32'h00000000;
      1356: value <= 32'h00000000;
      1357: value <= 32'h00000000;
      1358: value <= 32'h00000000;
      1359: value <= 32'h00000000;
      1360: value <= 32'h00000000;
      1361: value <= 32'h00000000;
      1362: value <= 32'h00000000;
      1363: value <= 32'h00000000;
      1364: value <= 32'h00000000;
      1365: value <= 32'h00000000;
      1366: value <= 32'h00000000;
      1367: value <= 32'h00000000;
      1368: value <= 32'h00000000;
      1369: value <= 32'h00000000;
      1370: value <= 32'h00000000;
      1371: value <= 32'h00000000;
      1372: value <= 32'h00000000;
      1373: value <= 32'h00000000;
      1374: value <= 32'h00000000;
      1375: value <= 32'h00000000;
      1376: value <= 32'h00000000;
      1377: value <= 32'h00000000;
      1378: value <= 32'h00000000;
      1379: value <= 32'h00000000;
      1380: value <= 32'h00000000;
      1381: value <= 32'h00000000;
      1382: value <= 32'h00000000;
      1383: value <= 32'h00000000;
      1384: value <= 32'h00000000;
      1385: value <= 32'h00000000;
      1386: value <= 32'h00000000;
      1387: value <= 32'h00000000;
      1388: value <= 32'h00000000;
      1389: value <= 32'h00000000;
      1390: value <= 32'h00000000;
      1391: value <= 32'h00000000;
      1392: value <= 32'h00000000;
      1393: value <= 32'h00000000;
      1394: value <= 32'h00000000;
      1395: value <= 32'h00000000;
      1396: value <= 32'h00000000;
      1397: value <= 32'h00000000;
      1398: value <= 32'h00000000;
      1399: value <= 32'h00000000;
      1400: value <= 32'h00000000;
      1401: value <= 32'h00000000;
      1402: value <= 32'h00000000;
      1403: value <= 32'h00000000;
      1404: value <= 32'h00000000;
      1405: value <= 32'h00000000;
      1406: value <= 32'h00000000;
      1407: value <= 32'h00000000;
      1408: value <= 32'h00000000;
      1409: value <= 32'h00000000;
      1410: value <= 32'h00000000;
      1411: value <= 32'h00000000;
      1412: value <= 32'h00000000;
      1413: value <= 32'h00000000;
      1414: value <= 32'h00000000;
      1415: value <= 32'h00000000;
      1416: value <= 32'h00000000;
      1417: value <= 32'h00000000;
      1418: value <= 32'h00000000;
      1419: value <= 32'h00000000;
      1420: value <= 32'h00000000;
      1421: value <= 32'h00000000;
      1422: value <= 32'h00000000;
      1423: value <= 32'h00000000;
      1424: value <= 32'h00000000;
      1425: value <= 32'h00000000;
      1426: value <= 32'h00000000;
      1427: value <= 32'h00000000;
      1428: value <= 32'h00000000;
      1429: value <= 32'h00000000;
      1430: value <= 32'h00000000;
      1431: value <= 32'h00000000;
      1432: value <= 32'h00000000;
      1433: value <= 32'h00000000;
      1434: value <= 32'h00000000;
      1435: value <= 32'h00000000;
      1436: value <= 32'h00000000;
      1437: value <= 32'h00000000;
      1438: value <= 32'h00000000;
      1439: value <= 32'h00000000;
      1440: value <= 32'h00000000;
      1441: value <= 32'h00000000;
      1442: value <= 32'h00000000;
      1443: value <= 32'h00000000;
      1444: value <= 32'h00000000;
      1445: value <= 32'h00000000;
      1446: value <= 32'h00000000;
      1447: value <= 32'h00000000;
      1448: value <= 32'h00000000;
      1449: value <= 32'h00000000;
      1450: value <= 32'h00000000;
      1451: value <= 32'h00000000;
      1452: value <= 32'h00000000;
      1453: value <= 32'h00000000;
      1454: value <= 32'h00000000;
      1455: value <= 32'h00000000;
      1456: value <= 32'h00000000;
      1457: value <= 32'h00000000;
      1458: value <= 32'h00000000;
      1459: value <= 32'h00000000;
      1460: value <= 32'h00000000;
      1461: value <= 32'h00000000;
      1462: value <= 32'h00000000;
      1463: value <= 32'h00000000;
      1464: value <= 32'h00000000;
      1465: value <= 32'h00000000;
      1466: value <= 32'h00000000;
      1467: value <= 32'h00000000;
      1468: value <= 32'h00000000;
      1469: value <= 32'h00000000;
      1470: value <= 32'h00000000;
      1471: value <= 32'h00000000;
      1472: value <= 32'h00000000;
      1473: value <= 32'h00000000;
      1474: value <= 32'h00000000;
      1475: value <= 32'h00000000;
      1476: value <= 32'h00000000;
      1477: value <= 32'h00000000;
      1478: value <= 32'h00000000;
      1479: value <= 32'h00000000;
      1480: value <= 32'h00000000;
      1481: value <= 32'h00000000;
      1482: value <= 32'h00000000;
      1483: value <= 32'h00000000;
      1484: value <= 32'h00000000;
      1485: value <= 32'h00000000;
      1486: value <= 32'h00000000;
      1487: value <= 32'h00000000;
      1488: value <= 32'h00000000;
      1489: value <= 32'h00000000;
      1490: value <= 32'h00000000;
      1491: value <= 32'h00000000;
      1492: value <= 32'h00000000;
      1493: value <= 32'h00000000;
      1494: value <= 32'h00000000;
      1495: value <= 32'h00000000;
      1496: value <= 32'h00000000;
      1497: value <= 32'h00000000;
      1498: value <= 32'h00000000;
      1499: value <= 32'h00000000;
      1500: value <= 32'h00000000;
      1501: value <= 32'h00000000;
      1502: value <= 32'h00000000;
      1503: value <= 32'h00000000;
      1504: value <= 32'h00000000;
      1505: value <= 32'h00000000;
      1506: value <= 32'h00000000;
      1507: value <= 32'h00000000;
      1508: value <= 32'h00000000;
      1509: value <= 32'h00000000;
      1510: value <= 32'h00000000;
      1511: value <= 32'h00000000;
      1512: value <= 32'h00000000;
      1513: value <= 32'h00000000;
      1514: value <= 32'h00000000;
      1515: value <= 32'h00000000;
      1516: value <= 32'h00000000;
      1517: value <= 32'h00000000;
      1518: value <= 32'h00000000;
      1519: value <= 32'h00000000;
      1520: value <= 32'h00000000;
      1521: value <= 32'h00000000;
      1522: value <= 32'h00000000;
      1523: value <= 32'h00000000;
      1524: value <= 32'h00000000;
      1525: value <= 32'h00000000;
      1526: value <= 32'h00000000;
      1527: value <= 32'h00000000;
      1528: value <= 32'h00000000;
      1529: value <= 32'h00000000;
      1530: value <= 32'h00000000;
      1531: value <= 32'h00000000;
      1532: value <= 32'h00000000;
      1533: value <= 32'h00000000;
      1534: value <= 32'h00000000;
      1535: value <= 32'h00000000;
      1536: value <= 32'h00000000;
      1537: value <= 32'h00000000;
      1538: value <= 32'h00000000;
      1539: value <= 32'h00000000;
      1540: value <= 32'h00000000;
      1541: value <= 32'h00000000;
      1542: value <= 32'h00000000;
      1543: value <= 32'h00000000;
      1544: value <= 32'h00000000;
      1545: value <= 32'h00000000;
      1546: value <= 32'h00000000;
      1547: value <= 32'h00000000;
      1548: value <= 32'h00000000;
      1549: value <= 32'h00000000;
      1550: value <= 32'h00000000;
      1551: value <= 32'h00000000;
      1552: value <= 32'h00000000;
      1553: value <= 32'h00000000;
      1554: value <= 32'h00000000;
      1555: value <= 32'h00000000;
      1556: value <= 32'h00000000;
      1557: value <= 32'h00000000;
      1558: value <= 32'h00000000;
      1559: value <= 32'h00000000;
      1560: value <= 32'h00000000;
      1561: value <= 32'h00000000;
      1562: value <= 32'h00000000;
      1563: value <= 32'h00000000;
      1564: value <= 32'h00000000;
      1565: value <= 32'h00000000;
      1566: value <= 32'h00000000;
      1567: value <= 32'h00000000;
      1568: value <= 32'h00000000;
      1569: value <= 32'h00000000;
      1570: value <= 32'h00000000;
      1571: value <= 32'h00000000;
      1572: value <= 32'h00000000;
      1573: value <= 32'h00000000;
      1574: value <= 32'h00000000;
      1575: value <= 32'h00000000;
      1576: value <= 32'h00000000;
      1577: value <= 32'h00000000;
      1578: value <= 32'h00000000;
      1579: value <= 32'h00000000;
      1580: value <= 32'h00000000;
      1581: value <= 32'h00000000;
      1582: value <= 32'h00000000;
      1583: value <= 32'h00000000;
      1584: value <= 32'h00000000;
      1585: value <= 32'h00000000;
      1586: value <= 32'h00000000;
      1587: value <= 32'h00000000;
      1588: value <= 32'h00000000;
      1589: value <= 32'h00000000;
      1590: value <= 32'h00000000;
      1591: value <= 32'h00000000;
      1592: value <= 32'h00000000;
      1593: value <= 32'h00000000;
      1594: value <= 32'h00000000;
      1595: value <= 32'h00000000;
      1596: value <= 32'h00000000;
      1597: value <= 32'h00000000;
      1598: value <= 32'h00000000;
      1599: value <= 32'h00000000;
      1600: value <= 32'h00000000;
      1601: value <= 32'h00000000;
      1602: value <= 32'h00000000;
      1603: value <= 32'h00000000;
      1604: value <= 32'h00000000;
      1605: value <= 32'h00000000;
      1606: value <= 32'h00000000;
      1607: value <= 32'h00000000;
      1608: value <= 32'h00000000;
      1609: value <= 32'h00000000;
      1610: value <= 32'h00000000;
      1611: value <= 32'h00000000;
      1612: value <= 32'h00000000;
      1613: value <= 32'h00000000;
      1614: value <= 32'h00000000;
      1615: value <= 32'h00000000;
      1616: value <= 32'h00000000;
      1617: value <= 32'h00000000;
      1618: value <= 32'h00000000;
      1619: value <= 32'h00000000;
      1620: value <= 32'h00000000;
      1621: value <= 32'h00000000;
      1622: value <= 32'h00000000;
      1623: value <= 32'h00000000;
      1624: value <= 32'h00000000;
      1625: value <= 32'h00000000;
      1626: value <= 32'h00000000;
      1627: value <= 32'h00000000;
      1628: value <= 32'h00000000;
      1629: value <= 32'h00000000;
      1630: value <= 32'h00000000;
      1631: value <= 32'h00000000;
      1632: value <= 32'h00000000;
      1633: value <= 32'h00000000;
      1634: value <= 32'h00000000;
      1635: value <= 32'h00000000;
      1636: value <= 32'h00000000;
      1637: value <= 32'h00000000;
      1638: value <= 32'h00000000;
      1639: value <= 32'h00000000;
      1640: value <= 32'h00000000;
      1641: value <= 32'h00000000;
      1642: value <= 32'h00000000;
      1643: value <= 32'h00000000;
      1644: value <= 32'h00000000;
      1645: value <= 32'h00000000;
      1646: value <= 32'h00000000;
      1647: value <= 32'h00000000;
      1648: value <= 32'h00000000;
      1649: value <= 32'h00000000;
      1650: value <= 32'h00000000;
      1651: value <= 32'h00000000;
      1652: value <= 32'h00000000;
      1653: value <= 32'h00000000;
      1654: value <= 32'h00000000;
      1655: value <= 32'h00000000;
      1656: value <= 32'h00000000;
      1657: value <= 32'h00000000;
      1658: value <= 32'h00000000;
      1659: value <= 32'h00000000;
      1660: value <= 32'h00000000;
      1661: value <= 32'h00000000;
      1662: value <= 32'h00000000;
      1663: value <= 32'h00000000;
      1664: value <= 32'h00000000;
      1665: value <= 32'h00000000;
      1666: value <= 32'h00000000;
      1667: value <= 32'h00000000;
      1668: value <= 32'h00000000;
      1669: value <= 32'h00000000;
      1670: value <= 32'h00000000;
      1671: value <= 32'h00000000;
      1672: value <= 32'h00000000;
      1673: value <= 32'h00000000;
      1674: value <= 32'h00000000;
      1675: value <= 32'h00000000;
      1676: value <= 32'h00000000;
      1677: value <= 32'h00000000;
      1678: value <= 32'h00000000;
      1679: value <= 32'h00000000;
      1680: value <= 32'h00000000;
      1681: value <= 32'h00000000;
      1682: value <= 32'h00000000;
      1683: value <= 32'h00000000;
      1684: value <= 32'h00000000;
      1685: value <= 32'h00000000;
      1686: value <= 32'h00000000;
      1687: value <= 32'h00000000;
      1688: value <= 32'h00000000;
      1689: value <= 32'h00000000;
      1690: value <= 32'h00000000;
      1691: value <= 32'h00000000;
      1692: value <= 32'h00000000;
      1693: value <= 32'h00000000;
      1694: value <= 32'h00000000;
      1695: value <= 32'h00000000;
      1696: value <= 32'h00000000;
      1697: value <= 32'h00000000;
      1698: value <= 32'h00000000;
      1699: value <= 32'h00000000;
      1700: value <= 32'h00000000;
      1701: value <= 32'h00000000;
      1702: value <= 32'h00000000;
      1703: value <= 32'h00000000;
      1704: value <= 32'h00000000;
      1705: value <= 32'h00000000;
      1706: value <= 32'h00000000;
      1707: value <= 32'h00000000;
      1708: value <= 32'h00000000;
      1709: value <= 32'h00000000;
      1710: value <= 32'h00000000;
      1711: value <= 32'h00000000;
      1712: value <= 32'h00000000;
      1713: value <= 32'h00000000;
      1714: value <= 32'h00000000;
      1715: value <= 32'h00000000;
      1716: value <= 32'h00000000;
      1717: value <= 32'h00000000;
      1718: value <= 32'h00000000;
      1719: value <= 32'h00000000;
      1720: value <= 32'h00000000;
      1721: value <= 32'h00000000;
      1722: value <= 32'h00000000;
      1723: value <= 32'h00000000;
      1724: value <= 32'h00000000;
      1725: value <= 32'h00000000;
      1726: value <= 32'h00000000;
      1727: value <= 32'h00000000;
      1728: value <= 32'h00000000;
      1729: value <= 32'h00000000;
      1730: value <= 32'h00000000;
      1731: value <= 32'h00000000;
      1732: value <= 32'h00000000;
      1733: value <= 32'h00000000;
      1734: value <= 32'h00000000;
      1735: value <= 32'h00000000;
      1736: value <= 32'h00000000;
      1737: value <= 32'h00000000;
      1738: value <= 32'h00000000;
      1739: value <= 32'h00000000;
      1740: value <= 32'h00000000;
      1741: value <= 32'h00000000;
      1742: value <= 32'h00000000;
      1743: value <= 32'h00000000;
      1744: value <= 32'h00000000;
      1745: value <= 32'h00000000;
      1746: value <= 32'h00000000;
      1747: value <= 32'h00000000;
      1748: value <= 32'h00000000;
      1749: value <= 32'h00000000;
      1750: value <= 32'h00000000;
      1751: value <= 32'h00000000;
      1752: value <= 32'h00000000;
      1753: value <= 32'h00000000;
      1754: value <= 32'h00000000;
      1755: value <= 32'h00000000;
      1756: value <= 32'h00000000;
      1757: value <= 32'h00000000;
      1758: value <= 32'h00000000;
      1759: value <= 32'h00000000;
      1760: value <= 32'h00000000;
      1761: value <= 32'h00000000;
      1762: value <= 32'h00000000;
      1763: value <= 32'h00000000;
      1764: value <= 32'h00000000;
      1765: value <= 32'h00000000;
      1766: value <= 32'h00000000;
      1767: value <= 32'h00000000;
      1768: value <= 32'h00000000;
      1769: value <= 32'h00000000;
      1770: value <= 32'h00000000;
      1771: value <= 32'h00000000;
      1772: value <= 32'h00000000;
      1773: value <= 32'h00000000;
      1774: value <= 32'h00000000;
      1775: value <= 32'h00000000;
      1776: value <= 32'h00000000;
      1777: value <= 32'h00000000;
      1778: value <= 32'h00000000;
      1779: value <= 32'h00000000;
      1780: value <= 32'h00000000;
      1781: value <= 32'h00000000;
      1782: value <= 32'h00000000;
      1783: value <= 32'h00000000;
      1784: value <= 32'h00000000;
      1785: value <= 32'h00000000;
      1786: value <= 32'h00000000;
      1787: value <= 32'h00000000;
      1788: value <= 32'h00000000;
      1789: value <= 32'h00000000;
      1790: value <= 32'h00000000;
      1791: value <= 32'h00000000;
      1792: value <= 32'h00000000;
      1793: value <= 32'h00000000;
      1794: value <= 32'h00000000;
      1795: value <= 32'h00000000;
      1796: value <= 32'h00000000;
      1797: value <= 32'h00000000;
      1798: value <= 32'h00000000;
      1799: value <= 32'h00000000;
      1800: value <= 32'h00000000;
      1801: value <= 32'h00000000;
      1802: value <= 32'h00000000;
      1803: value <= 32'h00000000;
      1804: value <= 32'h00000000;
      1805: value <= 32'h00000000;
      1806: value <= 32'h00000000;
      1807: value <= 32'h00000000;
      1808: value <= 32'h00000000;
      1809: value <= 32'h00000000;
      1810: value <= 32'h00000000;
      1811: value <= 32'h00000000;
      1812: value <= 32'h00000000;
      1813: value <= 32'h00000000;
      1814: value <= 32'h00000000;
      1815: value <= 32'h00000000;
      1816: value <= 32'h00000000;
      1817: value <= 32'h00000000;
      1818: value <= 32'h00000000;
      1819: value <= 32'h00000000;
      1820: value <= 32'h00000000;
      1821: value <= 32'h00000000;
      1822: value <= 32'h00000000;
      1823: value <= 32'h00000000;
      1824: value <= 32'h00000000;
      1825: value <= 32'h00000000;
      1826: value <= 32'h00000000;
      1827: value <= 32'h00000000;
      1828: value <= 32'h00000000;
      1829: value <= 32'h00000000;
      1830: value <= 32'h00000000;
      1831: value <= 32'h00000000;
      1832: value <= 32'h00000000;
      1833: value <= 32'h00000000;
      1834: value <= 32'h00000000;
      1835: value <= 32'h00000000;
      1836: value <= 32'h00000000;
      1837: value <= 32'h00000000;
      1838: value <= 32'h00000000;
      1839: value <= 32'h00000000;
      1840: value <= 32'h00000000;
      1841: value <= 32'h00000000;
      1842: value <= 32'h00000000;
      1843: value <= 32'h00000000;
      1844: value <= 32'h00000000;
      1845: value <= 32'h00000000;
      1846: value <= 32'h00000000;
      1847: value <= 32'h00000000;
      1848: value <= 32'h00000000;
      1849: value <= 32'h00000000;
      1850: value <= 32'h00000000;
      1851: value <= 32'h00000000;
      1852: value <= 32'h00000000;
      1853: value <= 32'h00000000;
      1854: value <= 32'h00000000;
      1855: value <= 32'h00000000;
      1856: value <= 32'h00000000;
      1857: value <= 32'h00000000;
      1858: value <= 32'h00000000;
      1859: value <= 32'h00000000;
      1860: value <= 32'h00000000;
      1861: value <= 32'h00000000;
      1862: value <= 32'h00000000;
      1863: value <= 32'h00000000;
      1864: value <= 32'h00000000;
      1865: value <= 32'h00000000;
      1866: value <= 32'h00000000;
      1867: value <= 32'h00000000;
      1868: value <= 32'h00000000;
      1869: value <= 32'h00000000;
      1870: value <= 32'h00000000;
      1871: value <= 32'h00000000;
      1872: value <= 32'h00000000;
      1873: value <= 32'h00000000;
      1874: value <= 32'h00000000;
      1875: value <= 32'h00000000;
      1876: value <= 32'h00000000;
      1877: value <= 32'h00000000;
      1878: value <= 32'h00000000;
      1879: value <= 32'h00000000;
      1880: value <= 32'h00000000;
      1881: value <= 32'h00000000;
      1882: value <= 32'h00000000;
      1883: value <= 32'h00000000;
      1884: value <= 32'h00000000;
      1885: value <= 32'h00000000;
      1886: value <= 32'h00000000;
      1887: value <= 32'h00000000;
      1888: value <= 32'h00000000;
      1889: value <= 32'h00000000;
      1890: value <= 32'h00000000;
      1891: value <= 32'h00000000;
      1892: value <= 32'h00000000;
      1893: value <= 32'h00000000;
      1894: value <= 32'h00000000;
      1895: value <= 32'h00000000;
      1896: value <= 32'h00000000;
      1897: value <= 32'h00000000;
      1898: value <= 32'h00000000;
      1899: value <= 32'h00000000;
      1900: value <= 32'h00000000;
      1901: value <= 32'h00000000;
      1902: value <= 32'h00000000;
      1903: value <= 32'h00000000;
      1904: value <= 32'h00000000;
      1905: value <= 32'h00000000;
      1906: value <= 32'h00000000;
      1907: value <= 32'h00000000;
      1908: value <= 32'h00000000;
      1909: value <= 32'h00000000;
      1910: value <= 32'h00000000;
      1911: value <= 32'h00000000;
      1912: value <= 32'h00000000;
      1913: value <= 32'h00000000;
      1914: value <= 32'h00000000;
      1915: value <= 32'h00000000;
      1916: value <= 32'h00000000;
      1917: value <= 32'h00000000;
      1918: value <= 32'h00000000;
      1919: value <= 32'h00000000;
      1920: value <= 32'h00000000;
      1921: value <= 32'h00000000;
      1922: value <= 32'h00000000;
      1923: value <= 32'h00000000;
      1924: value <= 32'h00000000;
      1925: value <= 32'h00000000;
      1926: value <= 32'h00000000;
      1927: value <= 32'h00000000;
      1928: value <= 32'h00000000;
      1929: value <= 32'h00000000;
      1930: value <= 32'h00000000;
      1931: value <= 32'h00000000;
      1932: value <= 32'h00000000;
      1933: value <= 32'h00000000;
      1934: value <= 32'h00000000;
      1935: value <= 32'h00000000;
      1936: value <= 32'h00000000;
      1937: value <= 32'h00000000;
      1938: value <= 32'h00000000;
      1939: value <= 32'h00000000;
      1940: value <= 32'h00000000;
      1941: value <= 32'h00000000;
      1942: value <= 32'h00000000;
      1943: value <= 32'h00000000;
      1944: value <= 32'h00000000;
      1945: value <= 32'h00000000;
      1946: value <= 32'h00000000;
      1947: value <= 32'h00000000;
      1948: value <= 32'h00000000;
      1949: value <= 32'h00000000;
      1950: value <= 32'h00000000;
      1951: value <= 32'h00000000;
      1952: value <= 32'h00000000;
      1953: value <= 32'h00000000;
      1954: value <= 32'h00000000;
      1955: value <= 32'h00000000;
      1956: value <= 32'h00000000;
      1957: value <= 32'h00000000;
      1958: value <= 32'h00000000;
      1959: value <= 32'h00000000;
      1960: value <= 32'h00000000;
      1961: value <= 32'h00000000;
      1962: value <= 32'h00000000;
      1963: value <= 32'h00000000;
      1964: value <= 32'h00000000;
      1965: value <= 32'h00000000;
      1966: value <= 32'h00000000;
      1967: value <= 32'h00000000;
      1968: value <= 32'h00000000;
      1969: value <= 32'h00000000;
      1970: value <= 32'h00000000;
      1971: value <= 32'h00000000;
      1972: value <= 32'h00000000;
      1973: value <= 32'h00000000;
      1974: value <= 32'h00000000;
      1975: value <= 32'h00000000;
      1976: value <= 32'h00000000;
      1977: value <= 32'h00000000;
      1978: value <= 32'h00000000;
      1979: value <= 32'h00000000;
      1980: value <= 32'h00000000;
      1981: value <= 32'h00000000;
      1982: value <= 32'h00000000;
      1983: value <= 32'h00000000;
      1984: value <= 32'h00000000;
      1985: value <= 32'h00000000;
      1986: value <= 32'h00000000;
      1987: value <= 32'h00000000;
      1988: value <= 32'h00000000;
      1989: value <= 32'h00000000;
      1990: value <= 32'h00000000;
      1991: value <= 32'h00000000;
      1992: value <= 32'h00000000;
      1993: value <= 32'h00000000;
      1994: value <= 32'h00000000;
      1995: value <= 32'h00000000;
      1996: value <= 32'h00000000;
      1997: value <= 32'h00000000;
      1998: value <= 32'h00000000;
      1999: value <= 32'h00000000;
      2000: value <= 32'h00000000;
      2001: value <= 32'h00000000;
      2002: value <= 32'h00000000;
      2003: value <= 32'h00000000;
      2004: value <= 32'h00000000;
      2005: value <= 32'h00000000;
      2006: value <= 32'h00000000;
      2007: value <= 32'h00000000;
      2008: value <= 32'h00000000;
      2009: value <= 32'h00000000;
      2010: value <= 32'h00000000;
      2011: value <= 32'h00000000;
      2012: value <= 32'h00000000;
      2013: value <= 32'h00000000;
      2014: value <= 32'h00000000;
      2015: value <= 32'h00000000;
      2016: value <= 32'h00000000;
      2017: value <= 32'h00000000;
      2018: value <= 32'h00000000;
      2019: value <= 32'h00000000;
      2020: value <= 32'h00000000;
      2021: value <= 32'h00000000;
      2022: value <= 32'h00000000;
      2023: value <= 32'h00000000;
      2024: value <= 32'h00000000;
      2025: value <= 32'h00000000;
      2026: value <= 32'h00000000;
      2027: value <= 32'h00000000;
      2028: value <= 32'h00000000;
      2029: value <= 32'h00000000;
      2030: value <= 32'h00000000;
      2031: value <= 32'h00000000;
      2032: value <= 32'h00000000;
      2033: value <= 32'h00000000;
      2034: value <= 32'h00000000;
      2035: value <= 32'h00000000;
      2036: value <= 32'h00000000;
      2037: value <= 32'h00000000;
      2038: value <= 32'h00000000;
      2039: value <= 32'h00000000;
      2040: value <= 32'h00000000;
      2041: value <= 32'h00000000;
      2042: value <= 32'h00000000;
      2043: value <= 32'h00000000;
      2044: value <= 32'h00000000;
      2045: value <= 32'h00000000;
      2046: value <= 32'h00000000;
      2047: value <= 32'h00000000;
      2048: value <= 32'h00000000;
      2049: value <= 32'h00000000;
      2050: value <= 32'h00000000;
      default: value <= 0;
    endcase
  end
endmodule
