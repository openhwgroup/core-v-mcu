module myDesign_QL_eFPGA_ArcticPro2_32X32_GF_22_QL_eFPGA (  CLK0, CLK1, CLK2, CLK3, CLK4, CLK5, fpgaio_data_0_i, fpgaio_data_1_i, fpgaio_data_2_i, fpgaio_data_3_i, fpgaio_data_4_i, fpgaio_data_5_i, fpgaio_data_6_i, fpgaio_data_7_i, udma_cfg_data_8_i, udma_cfg_data_9_i, udma_cfg_data_10_i, udma_cfg_data_11_i, udma_cfg_data_12_i, udma_cfg_data_13_i, udma_cfg_data_14_i, udma_cfg_data_15_i, udma_cfg_data_2_i, udma_cfg_data_3_i, udma_cfg_data_4_i, udma_cfg_data_5_i, udma_cfg_data_6_i, udma_cfg_data_7_i, udma_tx_lin_data_27_i, udma_tx_lin_data_28_i, udma_tx_lin_data_29_i, udma_tx_lin_data_30_i, udma_tx_lin_data_31_i, udma_rx_lin_ready_i, udma_cfg_data_0_i, udma_cfg_data_1_i, udma_tx_lin_data_21_i, udma_tx_lin_data_22_i, udma_tx_lin_data_23_i, udma_tx_lin_data_24_i, udma_tx_lin_data_25_i, udma_tx_lin_data_26_i, udma_tx_lin_data_13_i, udma_tx_lin_data_14_i, udma_tx_lin_data_15_i, udma_tx_lin_data_16_i, udma_tx_lin_data_17_i, udma_tx_lin_data_18_i, udma_tx_lin_data_19_i, udma_tx_lin_data_20_i, udma_tx_lin_data_7_i, udma_tx_lin_data_8_i, udma_tx_lin_data_9_i, udma_tx_lin_data_10_i, udma_tx_lin_data_11_i, udma_tx_lin_data_12_i, udma_tx_lin_valid_i, udma_tx_lin_data_0_i, udma_tx_lin_data_1_i, udma_tx_lin_data_2_i, udma_tx_lin_data_3_i, udma_tx_lin_data_4_i, udma_tx_lin_data_5_i, udma_tx_lin_data_6_i, apb_hwce_pwdata_0_i, apb_hwce_pwdata_1_i, apb_hwce_pwdata_2_i, apb_hwce_pwdata_3_i, apb_hwce_pwdata_4_i, apb_hwce_pwdata_5_i, apb_hwce_pwdata_6_i, apb_hwce_pwdata_7_i, apb_hwce_pwdata_8_i, apb_hwce_pwdata_9_i, apb_hwce_pwdata_10_i, apb_hwce_pwdata_11_i, apb_hwce_pwdata_12_i, apb_hwce_pwdata_13_i, apb_hwce_pwdata_14_i, apb_hwce_pwdata_15_i, apb_hwce_pwdata_16_i, apb_hwce_pwdata_17_i, apb_hwce_pwdata_18_i, apb_hwce_pwdata_19_i, apb_hwce_pwdata_20_i, apb_hwce_pwdata_21_i, apb_hwce_pwdata_22_i, apb_hwce_pwdata_23_i, apb_hwce_pwdata_24_i, apb_hwce_pwdata_25_i, apb_hwce_pwdata_26_i, apb_hwce_pwdata_27_i, apb_hwce_pwdata_28_i, apb_hwce_pwdata_29_i, apb_hwce_pwdata_30_i, apb_hwce_pwdata_31_i, apb_hwce_addr_0_i, apb_hwce_addr_1_i, apb_hwce_addr_2_i, apb_hwce_addr_3_i, apb_hwce_addr_4_i, apb_hwce_addr_5_i, apb_hwce_addr_6_i, apb_hwce_enable_i, apb_hwce_psel_i, apb_hwce_pstrb_i, apb_hwce_pwrite_i, fpgaio_data_28_i, fpgaio_data_29_i, fpgaio_data_30_i, fpgaio_data_31_i, fpgaio_data_32_i, fpgaio_data_33_i, fpgaio_data_34_i, fpgaio_data_35_i, fpgaio_data_36_i, fpgaio_data_37_i, fpgaio_data_38_i, fpgaio_data_39_i, fpgaio_data_40_i, fpgaio_data_41_i, fpgaio_data_42_i, RESET_LB, RESET_LT, fpgaio_data_20_i, fpgaio_data_21_i, fpgaio_data_22_i, fpgaio_data_23_i, fpgaio_data_24_i, fpgaio_data_25_i, fpgaio_data_26_i, fpgaio_data_27_i, udma_cfg_data_30_i, udma_cfg_data_31_i, fpgaio_data_16_i, fpgaio_data_17_i, fpgaio_data_18_i, fpgaio_data_19_i, udma_cfg_data_22_i, udma_cfg_data_23_i, udma_cfg_data_24_i, udma_cfg_data_25_i, udma_cfg_data_26_i, udma_cfg_data_27_i, udma_cfg_data_28_i, udma_cfg_data_29_i, udma_cfg_data_16_i, udma_cfg_data_17_i, udma_cfg_data_18_i, udma_cfg_data_19_i, udma_cfg_data_20_i, udma_cfg_data_21_i, tcdm_r_rdata_p3_8_i, tcdm_r_rdata_p3_9_i, tcdm_r_rdata_p3_10_i, tcdm_r_rdata_p3_11_i, tcdm_r_rdata_p3_12_i, tcdm_r_rdata_p3_13_i, tcdm_r_rdata_p3_14_i, tcdm_r_rdata_p3_15_i, tcdm_r_rdata_p3_2_i, tcdm_r_rdata_p3_3_i, tcdm_r_rdata_p3_4_i, tcdm_r_rdata_p3_5_i, tcdm_r_rdata_p3_6_i, tcdm_r_rdata_p3_7_i, tcdm_r_rdata_p2_28_i, tcdm_r_rdata_p2_29_i, tcdm_r_rdata_p2_30_i, tcdm_r_rdata_p2_31_i, tcdm_gnt_p2_i, tcdm_r_valid_p2_i, tcdm_r_rdata_p3_0_i, tcdm_r_rdata_p3_1_i, tcdm_r_rdata_p2_22_i, tcdm_r_rdata_p2_23_i, tcdm_r_rdata_p2_24_i, tcdm_r_rdata_p2_25_i, tcdm_r_rdata_p2_26_i, tcdm_r_rdata_p2_27_i, tcdm_r_rdata_p2_14_i, tcdm_r_rdata_p2_15_i, tcdm_r_rdata_p2_16_i, tcdm_r_rdata_p2_17_i, tcdm_r_rdata_p2_18_i, tcdm_r_rdata_p2_19_i, tcdm_r_rdata_p2_20_i, tcdm_r_rdata_p2_21_i, tcdm_r_rdata_p2_8_i, tcdm_r_rdata_p2_9_i, tcdm_r_rdata_p2_10_i, tcdm_r_rdata_p2_11_i, tcdm_r_rdata_p2_12_i, tcdm_r_rdata_p2_13_i, tcdm_r_rdata_p2_0_i, tcdm_r_rdata_p2_1_i, tcdm_r_rdata_p2_2_i, tcdm_r_rdata_p2_3_i, tcdm_r_rdata_p2_4_i, tcdm_r_rdata_p2_5_i, tcdm_r_rdata_p2_6_i, tcdm_r_rdata_p2_7_i, tcdm_r_rdata_p0_0_i, tcdm_r_rdata_p0_1_i, tcdm_r_rdata_p0_2_i, tcdm_r_rdata_p0_3_i, tcdm_r_rdata_p0_4_i, tcdm_r_rdata_p0_5_i, tcdm_r_rdata_p0_6_i, tcdm_r_rdata_p0_7_i, tcdm_r_rdata_p0_8_i, tcdm_r_rdata_p0_9_i, tcdm_r_rdata_p0_10_i, tcdm_r_rdata_p0_11_i, tcdm_r_rdata_p0_12_i, tcdm_r_rdata_p0_13_i, tcdm_r_rdata_p0_14_i, tcdm_r_rdata_p0_15_i, tcdm_r_rdata_p0_16_i, tcdm_r_rdata_p0_17_i, tcdm_r_rdata_p0_18_i, tcdm_r_rdata_p0_19_i, tcdm_r_rdata_p0_20_i, tcdm_r_rdata_p0_21_i, tcdm_r_rdata_p0_22_i, tcdm_r_rdata_p0_23_i, tcdm_r_rdata_p0_24_i, tcdm_r_rdata_p0_25_i, tcdm_r_rdata_p0_26_i, tcdm_r_rdata_p0_27_i, tcdm_r_rdata_p0_28_i, tcdm_r_rdata_p0_29_i, tcdm_r_rdata_p0_30_i, tcdm_r_rdata_p0_31_i, tcdm_gnt_p0_i, tcdm_r_valid_p0_i, tcdm_r_rdata_p1_0_i, tcdm_r_rdata_p1_1_i, tcdm_r_rdata_p1_2_i, tcdm_r_rdata_p1_3_i, tcdm_r_rdata_p1_4_i, tcdm_r_rdata_p1_5_i, tcdm_r_rdata_p1_6_i, tcdm_r_rdata_p1_7_i, tcdm_r_rdata_p1_8_i, tcdm_r_rdata_p1_9_i, tcdm_r_rdata_p1_10_i, tcdm_r_rdata_p1_11_i, tcdm_r_rdata_p1_12_i, tcdm_r_rdata_p1_13_i, tcdm_r_rdata_p1_14_i, tcdm_r_rdata_p1_15_i, tcdm_r_rdata_p1_16_i, tcdm_r_rdata_p1_17_i, tcdm_r_rdata_p1_18_i, tcdm_r_rdata_p1_19_i, tcdm_r_rdata_p1_20_i, tcdm_r_rdata_p1_21_i, tcdm_r_rdata_p1_22_i, tcdm_r_rdata_p1_23_i, tcdm_r_rdata_p1_24_i, tcdm_r_rdata_p1_25_i, tcdm_r_rdata_p1_26_i, tcdm_r_rdata_p1_27_i, tcdm_r_rdata_p1_28_i, tcdm_r_rdata_p1_29_i, tcdm_r_rdata_p1_30_i, tcdm_r_rdata_p1_31_i, tcdm_gnt_p1_i, tcdm_r_valid_p1_i, fpgaio_data_8_i, fpgaio_data_9_i, fpgaio_data_10_i, fpgaio_data_11_i, RESET_RB, fpgaio_data_14_i, fpgaio_data_15_i, RESET_RT, tcdm_r_rdata_p3_30_i, tcdm_r_rdata_p3_31_i, tcdm_gnt_p3_i, tcdm_r_valid_p3_i, fpgaio_data_12_i, fpgaio_data_13_i, tcdm_r_rdata_p3_22_i, tcdm_r_rdata_p3_23_i, tcdm_r_rdata_p3_24_i, tcdm_r_rdata_p3_25_i, tcdm_r_rdata_p3_26_i, tcdm_r_rdata_p3_27_i, tcdm_r_rdata_p3_28_i, tcdm_r_rdata_p3_29_i, tcdm_r_rdata_p3_16_i, tcdm_r_rdata_p3_17_i, tcdm_r_rdata_p3_18_i, tcdm_r_rdata_p3_19_i, tcdm_r_rdata_p3_20_i, tcdm_r_rdata_p3_21_i, MU0_MATHB_EFPGA_MAC_OUT_7_, MU0_MATHB_EFPGA_MAC_OUT_6_, MU0_MATHB_EFPGA_MAC_OUT_5_, MU0_MATHB_EFPGA_MAC_OUT_4_, MU0_MATHB_EFPGA_MAC_OUT_3_, MU0_MATHB_EFPGA_MAC_OUT_2_, MU0_MATHB_EFPGA_MAC_OUT_1_, MU0_MATHB_EFPGA_MAC_OUT_0_, MU0_TPRAM_EFPGA_COEF_R_DATA_31_, MU0_TPRAM_EFPGA_COEF_R_DATA_30_, MU0_TPRAM_EFPGA_COEF_R_DATA_29_, MU0_TPRAM_EFPGA_COEF_R_DATA_28_, MU0_TPRAM_EFPGA_COEF_R_DATA_27_, MU0_TPRAM_EFPGA_COEF_R_DATA_26_, MU0_TPRAM_EFPGA_COEF_R_DATA_25_, MU0_TPRAM_EFPGA_COEF_R_DATA_24_, MU0_TPRAM_EFPGA_COEF_R_DATA_23_, MU0_TPRAM_EFPGA_COEF_R_DATA_22_, MU0_TPRAM_EFPGA_COEF_R_DATA_21_, MU0_TPRAM_EFPGA_COEF_R_DATA_20_, MU0_TPRAM_EFPGA_COEF_R_DATA_19_, MU0_TPRAM_EFPGA_COEF_R_DATA_18_, MU0_TPRAM_EFPGA_COEF_R_DATA_17_, MU0_TPRAM_EFPGA_COEF_R_DATA_16_, MU0_TPRAM_EFPGA_COEF_R_DATA_15_, MU0_TPRAM_EFPGA_COEF_R_DATA_14_, MU0_TPRAM_EFPGA_COEF_R_DATA_13_, MU0_TPRAM_EFPGA_COEF_R_DATA_12_, MU0_TPRAM_EFPGA_COEF_R_DATA_11_, MU0_TPRAM_EFPGA_COEF_R_DATA_10_, MU0_TPRAM_EFPGA_COEF_R_DATA_9_, MU0_TPRAM_EFPGA_COEF_R_DATA_8_, MU0_TPRAM_EFPGA_COEF_R_DATA_7_, MU0_TPRAM_EFPGA_COEF_R_DATA_6_, MU0_TPRAM_EFPGA_COEF_R_DATA_5_, MU0_TPRAM_EFPGA_COEF_R_DATA_4_, MU0_TPRAM_EFPGA_COEF_R_DATA_3_, MU0_TPRAM_EFPGA_COEF_R_DATA_2_, MU0_TPRAM_EFPGA_COEF_R_DATA_1_, MU0_TPRAM_EFPGA_COEF_R_DATA_0_, MU1_TPRAM_EFPGA_OPER_R_DATA_31_, MU1_TPRAM_EFPGA_OPER_R_DATA_30_, MU1_TPRAM_EFPGA_OPER_R_DATA_29_, MU1_TPRAM_EFPGA_OPER_R_DATA_28_, MU1_TPRAM_EFPGA_OPER_R_DATA_27_, MU1_TPRAM_EFPGA_OPER_R_DATA_26_, MU1_TPRAM_EFPGA_OPER_R_DATA_25_, MU1_TPRAM_EFPGA_OPER_R_DATA_24_, MU1_TPRAM_EFPGA_OPER_R_DATA_23_, MU1_TPRAM_EFPGA_OPER_R_DATA_22_, MU1_TPRAM_EFPGA_OPER_R_DATA_21_, MU1_TPRAM_EFPGA_OPER_R_DATA_20_, MU1_TPRAM_EFPGA_OPER_R_DATA_19_, MU1_TPRAM_EFPGA_OPER_R_DATA_18_, MU1_TPRAM_EFPGA_OPER_R_DATA_17_, MU1_TPRAM_EFPGA_OPER_R_DATA_16_, MU1_TPRAM_EFPGA_OPER_R_DATA_15_, MU1_TPRAM_EFPGA_OPER_R_DATA_14_, MU1_TPRAM_EFPGA_OPER_R_DATA_13_, MU1_TPRAM_EFPGA_OPER_R_DATA_12_, MU0_TPRAM_EFPGA_OPER_R_DATA_31_, MU0_TPRAM_EFPGA_OPER_R_DATA_30_, MU0_TPRAM_EFPGA_OPER_R_DATA_29_, MU0_TPRAM_EFPGA_OPER_R_DATA_28_, MU1_TPRAM_EFPGA_OPER_R_DATA_11_, MU1_TPRAM_EFPGA_OPER_R_DATA_10_, MU1_TPRAM_EFPGA_OPER_R_DATA_9_, MU1_TPRAM_EFPGA_OPER_R_DATA_8_, MU1_TPRAM_EFPGA_OPER_R_DATA_7_, MU1_TPRAM_EFPGA_OPER_R_DATA_6_, MU1_TPRAM_EFPGA_OPER_R_DATA_5_, MU1_TPRAM_EFPGA_OPER_R_DATA_4_, MU1_TPRAM_EFPGA_OPER_R_DATA_3_, MU1_TPRAM_EFPGA_OPER_R_DATA_2_, MU1_TPRAM_EFPGA_OPER_R_DATA_1_, MU1_TPRAM_EFPGA_OPER_R_DATA_0_, MU1_MATHB_EFPGA_MAC_OUT_31_, MU1_MATHB_EFPGA_MAC_OUT_30_, MU1_MATHB_EFPGA_MAC_OUT_29_, MU1_MATHB_EFPGA_MAC_OUT_28_, MU1_MATHB_EFPGA_MAC_OUT_27_, MU1_MATHB_EFPGA_MAC_OUT_26_, MU1_MATHB_EFPGA_MAC_OUT_25_, MU1_MATHB_EFPGA_MAC_OUT_24_, MU1_MATHB_EFPGA_MAC_OUT_23_, MU1_MATHB_EFPGA_MAC_OUT_22_, MU1_MATHB_EFPGA_MAC_OUT_21_, MU1_MATHB_EFPGA_MAC_OUT_20_, MU1_MATHB_EFPGA_MAC_OUT_19_, MU1_MATHB_EFPGA_MAC_OUT_18_, MU1_MATHB_EFPGA_MAC_OUT_17_, MU1_MATHB_EFPGA_MAC_OUT_16_, MU1_MATHB_EFPGA_MAC_OUT_15_, MU1_MATHB_EFPGA_MAC_OUT_14_, MU1_MATHB_EFPGA_MAC_OUT_13_, MU1_MATHB_EFPGA_MAC_OUT_12_, MU1_MATHB_EFPGA_MAC_OUT_11_, MU1_MATHB_EFPGA_MAC_OUT_10_, MU1_MATHB_EFPGA_MAC_OUT_9_, MU1_MATHB_EFPGA_MAC_OUT_8_, MU1_MATHB_EFPGA_MAC_OUT_7_, MU1_MATHB_EFPGA_MAC_OUT_6_, MU1_MATHB_EFPGA_MAC_OUT_5_, MU1_MATHB_EFPGA_MAC_OUT_4_, MU1_MATHB_EFPGA_MAC_OUT_3_, MU1_MATHB_EFPGA_MAC_OUT_2_, MU1_MATHB_EFPGA_MAC_OUT_1_, MU1_MATHB_EFPGA_MAC_OUT_0_, MU1_TPRAM_EFPGA_COEF_R_DATA_31_, MU1_TPRAM_EFPGA_COEF_R_DATA_30_, MU1_TPRAM_EFPGA_COEF_R_DATA_29_, MU1_TPRAM_EFPGA_COEF_R_DATA_28_, MU1_TPRAM_EFPGA_COEF_R_DATA_27_, MU1_TPRAM_EFPGA_COEF_R_DATA_26_, MU1_TPRAM_EFPGA_COEF_R_DATA_25_, MU1_TPRAM_EFPGA_COEF_R_DATA_24_, MU1_TPRAM_EFPGA_COEF_R_DATA_23_, MU1_TPRAM_EFPGA_COEF_R_DATA_22_, MU1_TPRAM_EFPGA_COEF_R_DATA_21_, MU1_TPRAM_EFPGA_COEF_R_DATA_20_, MU1_TPRAM_EFPGA_COEF_R_DATA_19_, MU1_TPRAM_EFPGA_COEF_R_DATA_18_, MU0_TPRAM_EFPGA_OPER_R_DATA_27_, MU0_TPRAM_EFPGA_OPER_R_DATA_26_, MU0_TPRAM_EFPGA_OPER_R_DATA_25_, MU0_TPRAM_EFPGA_OPER_R_DATA_24_, MU0_TPRAM_EFPGA_OPER_R_DATA_23_, MU0_TPRAM_EFPGA_OPER_R_DATA_22_, MU0_TPRAM_EFPGA_OPER_R_DATA_21_, MU0_TPRAM_EFPGA_OPER_R_DATA_20_, MU1_TPRAM_EFPGA_COEF_R_DATA_17_, MU1_TPRAM_EFPGA_COEF_R_DATA_16_, MU1_TPRAM_EFPGA_COEF_R_DATA_15_, MU1_TPRAM_EFPGA_COEF_R_DATA_14_, MU1_TPRAM_EFPGA_COEF_R_DATA_13_, MU1_TPRAM_EFPGA_COEF_R_DATA_12_, MU1_TPRAM_EFPGA_COEF_R_DATA_11_, MU1_TPRAM_EFPGA_COEF_R_DATA_10_, MU1_TPRAM_EFPGA_COEF_R_DATA_9_, MU1_TPRAM_EFPGA_COEF_R_DATA_8_, MU1_TPRAM_EFPGA_COEF_R_DATA_7_, MU1_TPRAM_EFPGA_COEF_R_DATA_6_, MU1_TPRAM_EFPGA_COEF_R_DATA_5_, MU1_TPRAM_EFPGA_COEF_R_DATA_4_, MU1_TPRAM_EFPGA_COEF_R_DATA_3_, MU1_TPRAM_EFPGA_COEF_R_DATA_2_, MU1_TPRAM_EFPGA_COEF_R_DATA_1_, MU1_TPRAM_EFPGA_COEF_R_DATA_0_, MU0_TPRAM_EFPGA_OPER_R_DATA_19_, MU0_TPRAM_EFPGA_OPER_R_DATA_18_, MU0_TPRAM_EFPGA_OPER_R_DATA_17_, MU0_TPRAM_EFPGA_OPER_R_DATA_16_, MU0_TPRAM_EFPGA_OPER_R_DATA_15_, MU0_TPRAM_EFPGA_OPER_R_DATA_14_, MU0_TPRAM_EFPGA_OPER_R_DATA_13_, MU0_TPRAM_EFPGA_OPER_R_DATA_12_, MU0_TPRAM_EFPGA_OPER_R_DATA_11_, MU0_TPRAM_EFPGA_OPER_R_DATA_10_, MU0_TPRAM_EFPGA_OPER_R_DATA_9_, MU0_TPRAM_EFPGA_OPER_R_DATA_8_, MU0_TPRAM_EFPGA_OPER_R_DATA_7_, MU0_TPRAM_EFPGA_OPER_R_DATA_6_, MU0_TPRAM_EFPGA_OPER_R_DATA_5_, MU0_TPRAM_EFPGA_OPER_R_DATA_4_, MU0_TPRAM_EFPGA_OPER_R_DATA_3_, MU0_TPRAM_EFPGA_OPER_R_DATA_2_, MU0_TPRAM_EFPGA_OPER_R_DATA_1_, MU0_TPRAM_EFPGA_OPER_R_DATA_0_, MU0_MATHB_EFPGA_MAC_OUT_31_, MU0_MATHB_EFPGA_MAC_OUT_30_, MU0_MATHB_EFPGA_MAC_OUT_29_, MU0_MATHB_EFPGA_MAC_OUT_28_, MU0_MATHB_EFPGA_MAC_OUT_27_, MU0_MATHB_EFPGA_MAC_OUT_26_, MU0_MATHB_EFPGA_MAC_OUT_25_, MU0_MATHB_EFPGA_MAC_OUT_24_, MU0_MATHB_EFPGA_MAC_OUT_23_, MU0_MATHB_EFPGA_MAC_OUT_22_, MU0_MATHB_EFPGA_MAC_OUT_21_, MU0_MATHB_EFPGA_MAC_OUT_20_, MU0_MATHB_EFPGA_MAC_OUT_19_, MU0_MATHB_EFPGA_MAC_OUT_18_, MU0_MATHB_EFPGA_MAC_OUT_17_, MU0_MATHB_EFPGA_MAC_OUT_16_, MU0_MATHB_EFPGA_MAC_OUT_15_, MU0_MATHB_EFPGA_MAC_OUT_14_, MU0_MATHB_EFPGA_MAC_OUT_13_, MU0_MATHB_EFPGA_MAC_OUT_12_, MU0_MATHB_EFPGA_MAC_OUT_11_, MU0_MATHB_EFPGA_MAC_OUT_10_, MU0_MATHB_EFPGA_MAC_OUT_9_, MU0_MATHB_EFPGA_MAC_OUT_8_,  M_0_, BL_CLK, BL_DIN_0_, BL_DIN_10_, BL_DIN_11_, BL_DIN_12_, BL_DIN_13_, BL_DIN_14_, BL_DIN_15_, BL_DIN_16_, BL_DIN_17_, BL_DIN_18_, BL_DIN_19_, BL_DIN_1_, BL_DIN_20_, BL_DIN_21_, BL_DIN_22_, BL_DIN_23_, BL_DIN_24_, BL_DIN_25_, BL_DIN_26_, BL_DIN_27_, BL_DIN_28_, BL_DIN_29_, BL_DIN_2_, BL_DIN_30_, BL_DIN_31_, BL_DIN_3_, BL_DIN_4_, BL_DIN_5_, BL_DIN_6_, BL_DIN_7_, BL_DIN_8_, BL_DIN_9_, BL_PWRGATE_0_, BL_PWRGATE_1_, BL_PWRGATE_2_, BL_PWRGATE_3_, CLOAD_DIN_SEL, DIN_INT_L_ONLY, DIN_INT_R_ONLY, DIN_SLC_TB_INT, FB_CFG_DONE, FB_ISO_ENB, FB_SPE_IN_0_, FB_SPE_IN_1_, FB_SPE_IN_2_, FB_SPE_IN_3_, ISO_EN_0_, ISO_EN_1_, ISO_EN_2_, ISO_EN_3_, MLATCH, M_1_, M_2_, M_3_, M_4_, M_5_, NB, PB, PCHG_B, PI_PWR_0_, PI_PWR_1_, PI_PWR_2_, PI_PWR_3_, POR, PROG_0_, PROG_1_, PROG_2_, PROG_3_, PROG_IFX, PWR_GATE, RE, STM, VLP_CLKDIS_0_, VLP_CLKDIS_1_, VLP_CLKDIS_2_, VLP_CLKDIS_3_, VLP_CLKDIS_IFX, VLP_PWRDIS_0_, VLP_PWRDIS_1_, VLP_PWRDIS_2_, VLP_PWRDIS_3_, VLP_PWRDIS_IFX, VLP_SRDIS_0_, VLP_SRDIS_1_, VLP_SRDIS_2_, VLP_SRDIS_3_, VLP_SRDIS_IFX, WE, WE_INT, WL_CLK, WL_CLOAD_SEL_0_, WL_CLOAD_SEL_1_, WL_CLOAD_SEL_2_, WL_DIN_0_, WL_DIN_1_, WL_DIN_2_, WL_DIN_3_, WL_DIN_4_, WL_DIN_5_, WL_EN, WL_INT_DIN_SEL, WL_PWRGATE_0_, WL_PWRGATE_1_, WL_RESETB, WL_SEL_0_, WL_SEL_1_, WL_SEL_2_, WL_SEL_3_, WL_SEL_TB_INT, fpgaio_oe_0_o, fpgaio_data_0_o, fpgaio_oe_1_o, fpgaio_data_1_o, fpgaio_oe_2_o, fpgaio_data_2_o, fpgaio_oe_3_o, fpgaio_data_3_o, fpgaio_oe_4_o, fpgaio_data_4_o, fpgaio_oe_5_o, fpgaio_data_5_o, fpgaio_oe_6_o, fpgaio_data_6_o, fpgaio_oe_7_o, fpgaio_data_7_o, fpgaio_oe_20_o, fpgaio_data_20_o, fpgaio_oe_25_o, fpgaio_data_25_o, fpgaio_oe_26_o, fpgaio_data_26_o, fpgaio_oe_27_o, fpgaio_data_27_o, fpgaio_oe_21_o, fpgaio_data_21_o, fpgaio_oe_22_o, fpgaio_data_22_o, fpgaio_oe_23_o, fpgaio_data_23_o, fpgaio_oe_24_o, fpgaio_data_24_o, events_12_o, events_13_o, fpgaio_oe_19_o, fpgaio_data_19_o, events_14_o, events_15_o, fpgaio_oe_16_o, fpgaio_data_16_o, fpgaio_oe_17_o, fpgaio_data_17_o, fpgaio_oe_18_o, fpgaio_data_18_o, udma_cfg_data_26_o, udma_cfg_data_27_o, events_4_o, events_5_o, events_6_o, events_7_o, events_8_o, events_9_o, events_10_o, events_11_o, udma_cfg_data_28_o, udma_cfg_data_29_o, udma_cfg_data_30_o, udma_cfg_data_31_o, events_0_o, events_1_o, events_2_o, events_3_o, udma_cfg_data_14_o, udma_cfg_data_15_o, udma_cfg_data_24_o, udma_cfg_data_25_o, udma_cfg_data_16_o, udma_cfg_data_17_o, udma_cfg_data_18_o, udma_cfg_data_19_o, udma_cfg_data_20_o, udma_cfg_data_21_o, udma_cfg_data_22_o, udma_cfg_data_23_o, udma_rx_lin_data_28_o, udma_rx_lin_data_29_o, udma_cfg_data_6_o, udma_cfg_data_7_o, udma_cfg_data_8_o, udma_cfg_data_9_o, udma_cfg_data_10_o, udma_cfg_data_11_o, udma_cfg_data_12_o, udma_cfg_data_13_o, udma_rx_lin_data_30_o, udma_rx_lin_data_31_o, udma_cfg_data_0_o, udma_cfg_data_1_o, udma_cfg_data_2_o, udma_cfg_data_3_o, udma_cfg_data_4_o, udma_cfg_data_5_o, udma_rx_lin_data_16_o, udma_rx_lin_data_17_o, udma_rx_lin_data_26_o, udma_rx_lin_data_27_o, udma_rx_lin_data_18_o, udma_rx_lin_data_19_o, udma_rx_lin_data_20_o, udma_rx_lin_data_21_o, udma_rx_lin_data_22_o, udma_rx_lin_data_23_o, udma_rx_lin_data_24_o, udma_rx_lin_data_25_o, udma_tx_lin_ready_o, udma_rx_lin_valid_o, udma_rx_lin_data_8_o, udma_rx_lin_data_9_o, udma_rx_lin_data_10_o, udma_rx_lin_data_11_o, udma_rx_lin_data_12_o, udma_rx_lin_data_13_o, udma_rx_lin_data_14_o, udma_rx_lin_data_15_o, udma_rx_lin_data_0_o, udma_rx_lin_data_1_o, udma_rx_lin_data_2_o, udma_rx_lin_data_3_o, udma_rx_lin_data_4_o, udma_rx_lin_data_5_o, udma_rx_lin_data_6_o, udma_rx_lin_data_7_o, apb_hwce_prdata_0_o, apb_hwce_prdata_1_o, apb_hwce_prdata_10_o, apb_hwce_prdata_11_o, apb_hwce_prdata_2_o, apb_hwce_prdata_3_o, apb_hwce_prdata_4_o, apb_hwce_prdata_5_o, apb_hwce_prdata_6_o, apb_hwce_prdata_7_o, apb_hwce_prdata_8_o, apb_hwce_prdata_9_o, apb_hwce_prdata_12_o, apb_hwce_prdata_13_o, apb_hwce_prdata_22_o, apb_hwce_prdata_23_o, apb_hwce_prdata_24_o, apb_hwce_prdata_25_o, apb_hwce_prdata_26_o, apb_hwce_prdata_27_o, apb_hwce_prdata_28_o, apb_hwce_prdata_29_o, apb_hwce_prdata_14_o, apb_hwce_prdata_15_o, apb_hwce_prdata_16_o, apb_hwce_prdata_17_o, apb_hwce_prdata_18_o, apb_hwce_prdata_19_o, apb_hwce_prdata_20_o, apb_hwce_prdata_21_o, apb_hwce_prdata_30_o, apb_hwce_prdata_31_o, fpgaio_oe_31_o, fpgaio_data_31_o, apb_hwce_ready_o, apb_hwce_pslverr_o, fpgaio_oe_28_o, fpgaio_data_28_o, fpgaio_oe_29_o, fpgaio_data_29_o, fpgaio_oe_30_o, fpgaio_data_30_o, fpgaio_oe_32_o, fpgaio_data_32_o, fpgaio_oe_37_o, fpgaio_data_37_o, fpgaio_oe_38_o, fpgaio_data_38_o, fpgaio_oe_39_o, fpgaio_data_39_o, fpgaio_oe_40_o, fpgaio_data_40_o, fpgaio_oe_33_o, fpgaio_data_33_o, fpgaio_oe_34_o, fpgaio_data_34_o, fpgaio_oe_35_o, fpgaio_data_35_o, fpgaio_oe_36_o, fpgaio_data_36_o, fpgaio_oe_41_o, fpgaio_data_41_o, fpgaio_oe_42_o, fpgaio_data_42_o, tcdm_addr_p3_16_o, tcdm_wdata_p3_16_o, tcdm_wdata_p3_22_o, tcdm_wdata_p3_23_o, tcdm_wdata_p3_24_o, tcdm_wdata_p3_25_o, tcdm_wdata_p3_26_o, tcdm_wdata_p3_27_o, tcdm_wdata_p3_28_o, tcdm_wdata_p3_29_o, tcdm_addr_p3_17_o, tcdm_wdata_p3_17_o, tcdm_addr_p3_18_o, tcdm_wdata_p3_18_o, tcdm_addr_p3_19_o, tcdm_wdata_p3_19_o, tcdm_wdata_p3_20_o, tcdm_wdata_p3_21_o, tcdm_addr_p3_10_o, tcdm_wdata_p3_10_o, tcdm_addr_p3_15_o, tcdm_wdata_p3_15_o, tcdm_addr_p3_11_o, tcdm_wdata_p3_11_o, tcdm_addr_p3_12_o, tcdm_wdata_p3_12_o, tcdm_addr_p3_13_o, tcdm_wdata_p3_13_o, tcdm_addr_p3_14_o, tcdm_wdata_p3_14_o, tcdm_addr_p3_1_o, tcdm_wdata_p3_1_o, tcdm_addr_p3_6_o, tcdm_wdata_p3_6_o, tcdm_addr_p3_7_o, tcdm_wdata_p3_7_o, tcdm_addr_p3_8_o, tcdm_wdata_p3_8_o, tcdm_addr_p3_9_o, tcdm_wdata_p3_9_o, tcdm_addr_p3_2_o, tcdm_wdata_p3_2_o, tcdm_addr_p3_3_o, tcdm_wdata_p3_3_o, tcdm_addr_p3_4_o, tcdm_wdata_p3_4_o, tcdm_addr_p3_5_o, tcdm_wdata_p3_5_o, tcdm_wdata_p2_28_o, tcdm_wdata_p2_29_o, tcdm_addr_p3_0_o, tcdm_wdata_p3_0_o, tcdm_wdata_p2_30_o, tcdm_wdata_p2_31_o, tcdm_req_p2_o, tcdm_wen_p2_o, tcdm_be_p2_0_o, tcdm_be_p2_1_o, tcdm_be_p2_2_o, tcdm_be_p2_3_o, tcdm_addr_p2_15_o, tcdm_wdata_p2_15_o, tcdm_wdata_p2_20_o, tcdm_wdata_p2_21_o, tcdm_wdata_p2_22_o, tcdm_wdata_p2_23_o, tcdm_wdata_p2_24_o, tcdm_wdata_p2_25_o, tcdm_wdata_p2_26_o, tcdm_wdata_p2_27_o, tcdm_addr_p2_16_o, tcdm_wdata_p2_16_o, tcdm_addr_p2_17_o, tcdm_wdata_p2_17_o, tcdm_addr_p2_18_o, tcdm_wdata_p2_18_o, tcdm_addr_p2_19_o, tcdm_wdata_p2_19_o, tcdm_addr_p2_9_o, tcdm_wdata_p2_9_o, tcdm_addr_p2_14_o, tcdm_wdata_p2_14_o, tcdm_addr_p2_10_o, tcdm_wdata_p2_10_o, tcdm_addr_p2_11_o, tcdm_wdata_p2_11_o, tcdm_addr_p2_12_o, tcdm_wdata_p2_12_o, tcdm_addr_p2_13_o, tcdm_wdata_p2_13_o, tcdm_addr_p2_0_o, tcdm_wdata_p2_0_o, tcdm_addr_p2_5_o, tcdm_wdata_p2_5_o, tcdm_addr_p2_6_o, tcdm_wdata_p2_6_o, tcdm_addr_p2_7_o, tcdm_wdata_p2_7_o, tcdm_addr_p2_8_o, tcdm_wdata_p2_8_o, tcdm_addr_p2_1_o, tcdm_wdata_p2_1_o, tcdm_addr_p2_2_o, tcdm_wdata_p2_2_o, tcdm_addr_p2_3_o, tcdm_wdata_p2_3_o, tcdm_addr_p2_4_o, tcdm_wdata_p2_4_o, tcdm_addr_p0_0_o, tcdm_wdata_p0_0_o, tcdm_addr_p0_5_o, tcdm_wdata_p0_5_o, tcdm_addr_p0_1_o, tcdm_wdata_p0_1_o, tcdm_addr_p0_2_o, tcdm_wdata_p0_2_o, tcdm_addr_p0_3_o, tcdm_wdata_p0_3_o, tcdm_addr_p0_4_o, tcdm_wdata_p0_4_o, tcdm_addr_p0_6_o, tcdm_wdata_p0_6_o, tcdm_addr_p0_11_o, tcdm_wdata_p0_11_o, tcdm_addr_p0_12_o, tcdm_wdata_p0_12_o, tcdm_addr_p0_13_o, tcdm_wdata_p0_13_o, tcdm_addr_p0_14_o, tcdm_wdata_p0_14_o, tcdm_addr_p0_7_o, tcdm_wdata_p0_7_o, tcdm_addr_p0_8_o, tcdm_wdata_p0_8_o, tcdm_addr_p0_9_o, tcdm_wdata_p0_9_o, tcdm_addr_p0_10_o, tcdm_wdata_p0_10_o, tcdm_addr_p0_15_o, tcdm_wdata_p0_15_o, tcdm_wdata_p0_20_o, tcdm_wdata_p0_21_o, tcdm_addr_p0_16_o, tcdm_wdata_p0_16_o, tcdm_addr_p0_17_o, tcdm_wdata_p0_17_o, tcdm_addr_p0_18_o, tcdm_wdata_p0_18_o, tcdm_addr_p0_19_o, tcdm_wdata_p0_19_o, tcdm_wdata_p0_22_o, tcdm_wdata_p0_23_o, tcdm_req_p0_o, tcdm_wen_p0_o, tcdm_be_p0_0_o, tcdm_be_p0_1_o, tcdm_be_p0_2_o, tcdm_be_p0_3_o, tcdm_addr_p1_0_o, tcdm_wdata_p1_0_o, tcdm_wdata_p0_24_o, tcdm_wdata_p0_25_o, tcdm_wdata_p0_26_o, tcdm_wdata_p0_27_o, tcdm_wdata_p0_28_o, tcdm_wdata_p0_29_o, tcdm_wdata_p0_30_o, tcdm_wdata_p0_31_o, tcdm_addr_p1_1_o, tcdm_wdata_p1_1_o, tcdm_addr_p1_6_o, tcdm_wdata_p1_6_o, tcdm_addr_p1_2_o, tcdm_wdata_p1_2_o, tcdm_addr_p1_3_o, tcdm_wdata_p1_3_o, tcdm_addr_p1_4_o, tcdm_wdata_p1_4_o, tcdm_addr_p1_5_o, tcdm_wdata_p1_5_o, tcdm_addr_p1_7_o, tcdm_wdata_p1_7_o, tcdm_addr_p1_12_o, tcdm_wdata_p1_12_o, tcdm_addr_p1_13_o, tcdm_wdata_p1_13_o, tcdm_addr_p1_14_o, tcdm_wdata_p1_14_o, tcdm_addr_p1_15_o, tcdm_wdata_p1_15_o, tcdm_addr_p1_8_o, tcdm_wdata_p1_8_o, tcdm_addr_p1_9_o, tcdm_wdata_p1_9_o, tcdm_addr_p1_10_o, tcdm_wdata_p1_10_o, tcdm_addr_p1_11_o, tcdm_wdata_p1_11_o, tcdm_addr_p1_16_o, tcdm_wdata_p1_16_o, tcdm_wdata_p1_22_o, tcdm_wdata_p1_23_o, tcdm_addr_p1_17_o, tcdm_wdata_p1_17_o, tcdm_addr_p1_18_o, tcdm_wdata_p1_18_o, tcdm_addr_p1_19_o, tcdm_wdata_p1_19_o, tcdm_wdata_p1_20_o, tcdm_wdata_p1_21_o, tcdm_wdata_p1_24_o, tcdm_wdata_p1_25_o, tcdm_be_p1_0_o, tcdm_be_p1_1_o, tcdm_be_p1_2_o, tcdm_be_p1_3_o, fpgaio_oe_8_o, fpgaio_data_8_o, fpgaio_oe_9_o, fpgaio_data_9_o, tcdm_wdata_p1_26_o, tcdm_wdata_p1_27_o, tcdm_wdata_p1_28_o, tcdm_wdata_p1_29_o, tcdm_wdata_p1_30_o, tcdm_wdata_p1_31_o, tcdm_req_p1_o, tcdm_wen_p1_o, fpgaio_oe_10_o, fpgaio_data_10_o, fpgaio_oe_11_o, fpgaio_data_11_o, fpgaio_oe_14_o, fpgaio_data_14_o, fpgaio_oe_15_o, fpgaio_data_15_o, tcdm_wdata_p3_30_o, tcdm_wdata_p3_31_o, fpgaio_oe_13_o, fpgaio_data_13_o, tcdm_req_p3_o, tcdm_wen_p3_o, tcdm_be_p3_0_o, tcdm_be_p3_1_o, tcdm_be_p3_2_o, tcdm_be_p3_3_o, fpgaio_oe_12_o, fpgaio_data_12_o, MU0_EFPGA_MATHB_COEF_DATA_23_, MU0_EFPGA_MATHB_COEF_DATA_22_, MU0_EFPGA_MATHB_COEF_DATA_13_, MU0_EFPGA_MATHB_COEF_DATA_12_, MU0_EFPGA_MATHB_COEF_DATA_11_, MU0_EFPGA_MATHB_COEF_DATA_10_, MU0_EFPGA_MATHB_COEF_DATA_9_, MU0_EFPGA_MATHB_COEF_DATA_8_, MU0_EFPGA_MATHB_COEF_DATA_7_, MU0_EFPGA_MATHB_COEF_DATA_6_, MU0_EFPGA_MATHB_COEF_DATA_21_, MU0_EFPGA_MATHB_COEF_DATA_20_, MU0_EFPGA_MATHB_COEF_DATA_19_, MU0_EFPGA_MATHB_COEF_DATA_18_, MU0_EFPGA_MATHB_COEF_DATA_17_, MU0_EFPGA_MATHB_COEF_DATA_16_, MU0_EFPGA_MATHB_COEF_DATA_15_, MU0_EFPGA_MATHB_COEF_DATA_14_, MU0_EFPGA_MATHB_COEF_DATA_5_, MU0_EFPGA_MATHB_COEF_DATA_4_, MU0_EFPGA_TPRAM_COEF_W_DATA_31_, MU0_EFPGA_TPRAM_COEF_W_DATA_30_, MU0_EFPGA_MATHB_COEF_DATA_3_, MU0_EFPGA_MATHB_COEF_DATA_2_, MU0_EFPGA_MATHB_COEF_DATA_1_, MU0_EFPGA_MATHB_COEF_DATA_0_, MU0_EFPGA_MATHB_DATAOUT_SEL_1_, MU0_EFPGA_MATHB_DATAOUT_SEL_0_, MU0_EFPGA_TPRAM_COEF_W_MODE_1_, MU0_EFPGA_TPRAM_COEF_W_MODE_0_, MU0_EFPGA_TPRAM_COEF_W_DATA_29_, MU0_EFPGA_TPRAM_COEF_W_DATA_28_, MU0_EFPGA_TPRAM_COEF_W_DATA_19_, MU0_EFPGA_TPRAM_COEF_W_DATA_18_, MU0_EFPGA_TPRAM_COEF_W_DATA_17_, MU0_EFPGA_TPRAM_COEF_W_DATA_16_, MU0_EFPGA_TPRAM_COEF_W_DATA_15_, MU0_EFPGA_TPRAM_COEF_W_DATA_14_, MU0_EFPGA_TPRAM_COEF_W_DATA_13_, MU0_EFPGA_TPRAM_COEF_W_DATA_12_, MU0_EFPGA_TPRAM_COEF_W_DATA_27_, MU0_EFPGA_TPRAM_COEF_W_DATA_26_, MU0_EFPGA_TPRAM_COEF_W_DATA_25_, MU0_EFPGA_TPRAM_COEF_W_DATA_24_, MU0_EFPGA_TPRAM_COEF_W_DATA_23_, MU0_EFPGA_TPRAM_COEF_W_DATA_22_, MU0_EFPGA_TPRAM_COEF_W_DATA_21_, MU0_EFPGA_TPRAM_COEF_W_DATA_20_, MU0_EFPGA_TPRAM_COEF_W_DATA_11_, MU0_EFPGA_TPRAM_COEF_W_DATA_10_, MU0_EFPGA_TPRAM_COEF_W_DATA_1_, MU0_EFPGA_TPRAM_COEF_W_DATA_0_, MU0_EFPGA_TPRAM_COEF_W_DATA_9_, MU0_EFPGA_TPRAM_COEF_W_DATA_8_, MU0_EFPGA_TPRAM_COEF_W_DATA_7_, MU0_EFPGA_TPRAM_COEF_W_DATA_6_, MU0_EFPGA_TPRAM_COEF_W_DATA_5_, MU0_EFPGA_TPRAM_COEF_W_DATA_4_, MU0_EFPGA_TPRAM_COEF_W_DATA_3_, MU0_EFPGA_TPRAM_COEF_W_DATA_2_, MU0_EFPGA_TPRAM_COEF_W_CLK, MU0_EFPGA_TPRAM_COEF_W_ADDR_11_, MU0_EFPGA_TPRAM_COEF_W_ADDR_2_, MU0_EFPGA_TPRAM_COEF_W_ADDR_1_, MU0_EFPGA_TPRAM_COEF_W_ADDR_0_, MU0_EFPGA_TPRAM_COEF_WE, MU0_EFPGA_TPRAM_COEF_WDSEL, MU0_EFPGA_TPRAM_COEF_R_MODE_1_, MU0_EFPGA_TPRAM_COEF_R_MODE_0_, MU0_EFPGA_TPRAM_COEF_R_CLK, MU0_EFPGA_TPRAM_COEF_W_ADDR_10_, MU0_EFPGA_TPRAM_COEF_W_ADDR_9_, MU0_EFPGA_TPRAM_COEF_W_ADDR_8_, MU0_EFPGA_TPRAM_COEF_W_ADDR_7_, MU0_EFPGA_TPRAM_COEF_W_ADDR_6_, MU0_EFPGA_TPRAM_COEF_W_ADDR_5_, MU0_EFPGA_TPRAM_COEF_W_ADDR_4_, MU0_EFPGA_TPRAM_COEF_W_ADDR_3_, MU0_EFPGA_TPRAM_COEF_R_ADDR_11_, MU0_EFPGA_TPRAM_COEF_R_ADDR_10_, MU0_EFPGA_TPRAM_COEF_R_ADDR_1_, MU0_EFPGA_TPRAM_COEF_R_ADDR_0_, MU0_EFPGA_TPRAM_COEF_R_ADDR_9_, MU0_EFPGA_TPRAM_COEF_R_ADDR_8_, MU0_EFPGA_TPRAM_COEF_R_ADDR_7_, MU0_EFPGA_TPRAM_COEF_R_ADDR_6_, MU0_EFPGA_TPRAM_COEF_R_ADDR_5_, MU0_EFPGA_TPRAM_COEF_R_ADDR_4_, MU0_EFPGA_TPRAM_COEF_R_ADDR_3_, MU0_EFPGA_TPRAM_COEF_R_ADDR_2_, MU0_EFPGA_TPRAM_COEF_POWERDN, MU1_EFPGA_TPRAM_OPER_W_MODE_1_, MU1_EFPGA_TPRAM_OPER_W_MODE_0_, MU1_EFPGA_TPRAM_OPER_W_DATA_23_, MU1_EFPGA_TPRAM_OPER_W_DATA_22_, MU1_EFPGA_TPRAM_OPER_W_DATA_31_, MU1_EFPGA_TPRAM_OPER_W_DATA_30_, MU1_EFPGA_TPRAM_OPER_W_DATA_29_, MU1_EFPGA_TPRAM_OPER_W_DATA_28_, MU1_EFPGA_TPRAM_OPER_W_DATA_27_, MU1_EFPGA_TPRAM_OPER_W_DATA_26_, MU1_EFPGA_TPRAM_OPER_W_DATA_25_, MU1_EFPGA_TPRAM_OPER_W_DATA_24_, MU1_EFPGA_TPRAM_OPER_W_DATA_21_, MU1_EFPGA_TPRAM_OPER_W_DATA_20_, MU1_EFPGA_TPRAM_OPER_W_DATA_11_, MU1_EFPGA_TPRAM_OPER_W_DATA_10_, MU1_EFPGA_TPRAM_OPER_W_DATA_9_, MU1_EFPGA_TPRAM_OPER_W_DATA_8_, MU1_EFPGA_TPRAM_OPER_W_DATA_7_, MU1_EFPGA_TPRAM_OPER_W_DATA_6_, MU1_EFPGA_TPRAM_OPER_W_DATA_5_, MU1_EFPGA_TPRAM_OPER_W_DATA_4_, MU1_EFPGA_TPRAM_OPER_W_DATA_19_, MU1_EFPGA_TPRAM_OPER_W_DATA_18_, MU1_EFPGA_TPRAM_OPER_W_DATA_17_, MU1_EFPGA_TPRAM_OPER_W_DATA_16_, MU1_EFPGA_TPRAM_OPER_W_DATA_15_, MU1_EFPGA_TPRAM_OPER_W_DATA_14_, MU1_EFPGA_TPRAM_OPER_W_DATA_13_, MU1_EFPGA_TPRAM_OPER_W_DATA_12_, MU1_EFPGA_TPRAM_OPER_W_DATA_3_, MU1_EFPGA_TPRAM_OPER_W_DATA_2_, MU1_EFPGA_TPRAM_OPER_W_ADDR_6_, MU1_EFPGA_TPRAM_OPER_W_ADDR_5_, MU1_EFPGA_TPRAM_OPER_W_DATA_1_, MU1_EFPGA_TPRAM_OPER_W_DATA_0_, MU1_EFPGA_TPRAM_OPER_W_CLK, MU1_EFPGA_TPRAM_OPER_W_ADDR_11_, MU1_EFPGA_TPRAM_OPER_W_ADDR_10_, MU1_EFPGA_TPRAM_OPER_W_ADDR_9_, MU1_EFPGA_TPRAM_OPER_W_ADDR_8_, MU1_EFPGA_TPRAM_OPER_W_ADDR_7_, MU1_EFPGA_TPRAM_OPER_W_ADDR_4_, MU1_EFPGA_TPRAM_OPER_W_ADDR_3_, MU1_EFPGA_TPRAM_OPER_R_ADDR_11_, MU1_EFPGA_TPRAM_OPER_R_ADDR_10_, MU1_EFPGA_TPRAM_OPER_R_ADDR_9_, MU1_EFPGA_TPRAM_OPER_R_ADDR_8_, MU1_EFPGA_TPRAM_OPER_R_ADDR_7_, MU1_EFPGA_TPRAM_OPER_R_ADDR_6_, MU1_EFPGA_TPRAM_OPER_R_ADDR_5_, MU1_EFPGA_TPRAM_OPER_R_ADDR_4_, MU1_EFPGA_TPRAM_OPER_W_ADDR_2_, MU1_EFPGA_TPRAM_OPER_W_ADDR_1_, MU1_EFPGA_TPRAM_OPER_W_ADDR_0_, MU1_EFPGA_TPRAM_OPER_WE, MU1_EFPGA_TPRAM_OPER_WDSEL, MU1_EFPGA_TPRAM_OPER_R_MODE_1_, MU1_EFPGA_TPRAM_OPER_R_MODE_0_, MU1_EFPGA_TPRAM_OPER_R_CLK, MU1_EFPGA_TPRAM_OPER_R_ADDR_3_, MU1_EFPGA_TPRAM_OPER_R_ADDR_2_, MU1_EFPGA_MATHB_MAC_OUT_SEL_2_, MU1_EFPGA_MATHB_MAC_OUT_SEL_1_, MU1_EFPGA_TPRAM_OPER_R_ADDR_1_, MU1_EFPGA_TPRAM_OPER_R_ADDR_0_, MU1_EFPGA_TPRAM_OPER_POWERDN, MU1_EFPGA2MATHB_CLK, MU1_EFPGA_MATHB_CLK_EN, MU1_EFPGA_MATHB_MAC_OUT_SEL_5_, MU1_EFPGA_MATHB_MAC_OUT_SEL_4_, MU1_EFPGA_MATHB_MAC_OUT_SEL_3_, MU1_EFPGA_MATHB_MAC_OUT_SEL_0_, MU1_EFPGA_MATHB_MAC_ACC_SAT, MU1_EFPGA_MATHB_OPER_DATA_26_, MU1_EFPGA_MATHB_OPER_DATA_25_, MU1_EFPGA_MATHB_OPER_DATA_24_, MU1_EFPGA_MATHB_OPER_DATA_23_, MU1_EFPGA_MATHB_OPER_DATA_22_, MU1_EFPGA_MATHB_OPER_DATA_21_, MU1_EFPGA_MATHB_OPER_DATA_20_, MU1_EFPGA_MATHB_OPER_DATA_19_, MU1_EFPGA_MATHB_MAC_ACC_RND, MU1_EFPGA_MATHB_MAC_ACC_CLEAR, MU1_EFPGA_MATHB_OPER_SEL, MU1_EFPGA_MATHB_OPER_DATA_31_, MU1_EFPGA_MATHB_OPER_DATA_30_, MU1_EFPGA_MATHB_OPER_DATA_29_, MU1_EFPGA_MATHB_OPER_DATA_28_, MU1_EFPGA_MATHB_OPER_DATA_27_, MU1_EFPGA_MATHB_OPER_DATA_18_, MU1_EFPGA_MATHB_OPER_DATA_17_, MU1_EFPGA_MATHB_OPER_DATA_8_, MU1_EFPGA_MATHB_OPER_DATA_7_, MU1_EFPGA_MATHB_OPER_DATA_16_, MU1_EFPGA_MATHB_OPER_DATA_15_, MU1_EFPGA_MATHB_OPER_DATA_14_, MU1_EFPGA_MATHB_OPER_DATA_13_, MU1_EFPGA_MATHB_OPER_DATA_12_, MU1_EFPGA_MATHB_OPER_DATA_11_, MU1_EFPGA_MATHB_OPER_DATA_10_, MU1_EFPGA_MATHB_OPER_DATA_9_, MU1_EFPGA_MATHB_OPER_DATA_6_, MU1_EFPGA_MATHB_OPER_DATA_5_, MU1_EFPGA_MATHB_COEF_DATA_29_, MU1_EFPGA_MATHB_COEF_DATA_28_, MU1_EFPGA_MATHB_COEF_DATA_27_, MU1_EFPGA_MATHB_COEF_DATA_26_, MU1_EFPGA_MATHB_COEF_DATA_25_, MU1_EFPGA_MATHB_COEF_DATA_24_, MU1_EFPGA_MATHB_COEF_DATA_23_, MU1_EFPGA_MATHB_COEF_DATA_22_, MU1_EFPGA_MATHB_OPER_DATA_4_, MU1_EFPGA_MATHB_OPER_DATA_3_, MU1_EFPGA_MATHB_OPER_DATA_2_, MU1_EFPGA_MATHB_OPER_DATA_1_, MU1_EFPGA_MATHB_OPER_DATA_0_, MU1_EFPGA_MATHB_COEF_SEL, MU1_EFPGA_MATHB_COEF_DATA_31_, MU1_EFPGA_MATHB_COEF_DATA_30_, MU1_EFPGA_MATHB_COEF_DATA_21_, MU1_EFPGA_MATHB_COEF_DATA_20_, MU1_EFPGA_MATHB_COEF_DATA_11_, MU1_EFPGA_MATHB_COEF_DATA_10_, MU1_EFPGA_MATHB_COEF_DATA_19_, MU1_EFPGA_MATHB_COEF_DATA_18_, MU1_EFPGA_MATHB_COEF_DATA_17_, MU1_EFPGA_MATHB_COEF_DATA_16_, MU1_EFPGA_MATHB_COEF_DATA_15_, MU1_EFPGA_MATHB_COEF_DATA_14_, MU1_EFPGA_MATHB_COEF_DATA_13_, MU1_EFPGA_MATHB_COEF_DATA_12_, MU1_EFPGA_MATHB_COEF_DATA_9_, MU1_EFPGA_MATHB_COEF_DATA_8_, MU1_EFPGA_MATHB_DATAOUT_SEL_1_, MU1_EFPGA_MATHB_DATAOUT_SEL_0_, MU1_EFPGA_TPRAM_COEF_W_MODE_1_, MU1_EFPGA_TPRAM_COEF_W_MODE_0_, MU1_EFPGA_TPRAM_COEF_W_DATA_31_, MU1_EFPGA_TPRAM_COEF_W_DATA_30_, MU1_EFPGA_TPRAM_COEF_W_DATA_29_, MU1_EFPGA_TPRAM_COEF_W_DATA_28_, MU1_EFPGA_MATHB_COEF_DATA_7_, MU1_EFPGA_MATHB_COEF_DATA_6_, MU1_EFPGA_MATHB_COEF_DATA_5_, MU1_EFPGA_MATHB_COEF_DATA_4_, MU1_EFPGA_MATHB_COEF_DATA_3_, MU1_EFPGA_MATHB_COEF_DATA_2_, MU1_EFPGA_MATHB_COEF_DATA_1_, MU1_EFPGA_MATHB_COEF_DATA_0_, MU1_EFPGA_TPRAM_COEF_W_DATA_27_, MU1_EFPGA_TPRAM_COEF_W_DATA_26_, MU1_EFPGA_TPRAM_COEF_W_DATA_17_, MU1_EFPGA_TPRAM_COEF_W_DATA_16_, MU1_EFPGA_TPRAM_COEF_W_DATA_25_, MU1_EFPGA_TPRAM_COEF_W_DATA_24_, MU1_EFPGA_TPRAM_COEF_W_DATA_23_, MU1_EFPGA_TPRAM_COEF_W_DATA_22_, MU1_EFPGA_TPRAM_COEF_W_DATA_21_, MU1_EFPGA_TPRAM_COEF_W_DATA_20_, MU1_EFPGA_TPRAM_COEF_W_DATA_19_, MU1_EFPGA_TPRAM_COEF_W_DATA_18_, MU1_EFPGA_TPRAM_COEF_W_DATA_15_, MU1_EFPGA_TPRAM_COEF_W_DATA_14_, MU1_EFPGA_TPRAM_COEF_W_DATA_5_, MU1_EFPGA_TPRAM_COEF_W_DATA_4_, MU1_EFPGA_TPRAM_COEF_W_DATA_3_, MU1_EFPGA_TPRAM_COEF_W_DATA_2_, MU1_EFPGA_TPRAM_COEF_W_DATA_1_, MU1_EFPGA_TPRAM_COEF_W_DATA_0_, MU1_EFPGA_TPRAM_COEF_W_CLK, MU1_EFPGA_TPRAM_COEF_W_ADDR_11_, MU1_EFPGA_TPRAM_COEF_W_DATA_13_, MU1_EFPGA_TPRAM_COEF_W_DATA_12_, MU1_EFPGA_TPRAM_COEF_W_DATA_11_, MU1_EFPGA_TPRAM_COEF_W_DATA_10_, MU1_EFPGA_TPRAM_COEF_W_DATA_9_, MU1_EFPGA_TPRAM_COEF_W_DATA_8_, MU1_EFPGA_TPRAM_COEF_W_DATA_7_, MU1_EFPGA_TPRAM_COEF_W_DATA_6_, MU1_EFPGA_TPRAM_COEF_W_ADDR_10_, MU1_EFPGA_TPRAM_COEF_W_ADDR_9_, MU1_EFPGA_TPRAM_COEF_W_ADDR_0_, MU1_EFPGA_TPRAM_COEF_WE, MU1_EFPGA_TPRAM_COEF_W_ADDR_8_, MU1_EFPGA_TPRAM_COEF_W_ADDR_7_, MU1_EFPGA_TPRAM_COEF_W_ADDR_6_, MU1_EFPGA_TPRAM_COEF_W_ADDR_5_, MU1_EFPGA_TPRAM_COEF_W_ADDR_4_, MU1_EFPGA_TPRAM_COEF_W_ADDR_3_, MU1_EFPGA_TPRAM_COEF_W_ADDR_2_, MU1_EFPGA_TPRAM_COEF_W_ADDR_1_, MU0_EFPGA_TPRAM_OPER_W_DATA_25_, MU0_EFPGA_TPRAM_OPER_W_DATA_24_, MU0_EFPGA_TPRAM_OPER_W_DATA_23_, MU0_EFPGA_TPRAM_OPER_W_DATA_22_, MU0_EFPGA_TPRAM_OPER_W_DATA_21_, MU0_EFPGA_TPRAM_OPER_W_DATA_20_, MU0_EFPGA_TPRAM_OPER_W_DATA_19_, MU0_EFPGA_TPRAM_OPER_W_DATA_18_, MU0_EFPGA_TPRAM_OPER_W_MODE_1_, MU0_EFPGA_TPRAM_OPER_W_MODE_0_, MU0_EFPGA_TPRAM_OPER_W_DATA_31_, MU0_EFPGA_TPRAM_OPER_W_DATA_30_, MU0_EFPGA_TPRAM_OPER_W_DATA_29_, MU0_EFPGA_TPRAM_OPER_W_DATA_28_, MU0_EFPGA_TPRAM_OPER_W_DATA_27_, MU0_EFPGA_TPRAM_OPER_W_DATA_26_, MU1_EFPGA_TPRAM_COEF_WDSEL, MU1_EFPGA_TPRAM_COEF_R_MODE_1_, MU1_EFPGA_TPRAM_COEF_R_ADDR_5_, MU1_EFPGA_TPRAM_COEF_R_ADDR_4_, MU1_EFPGA_TPRAM_COEF_R_ADDR_3_, MU1_EFPGA_TPRAM_COEF_R_ADDR_2_, MU1_EFPGA_TPRAM_COEF_R_ADDR_1_, MU1_EFPGA_TPRAM_COEF_R_ADDR_0_, MU1_EFPGA_TPRAM_COEF_POWERDN, MU1_EFPGA_TPRAM_COEF_R_MODE_0_, MU1_EFPGA_TPRAM_COEF_R_CLK, MU1_EFPGA_TPRAM_COEF_R_ADDR_11_, MU1_EFPGA_TPRAM_COEF_R_ADDR_10_, MU1_EFPGA_TPRAM_COEF_R_ADDR_9_, MU1_EFPGA_TPRAM_COEF_R_ADDR_8_, MU1_EFPGA_TPRAM_COEF_R_ADDR_7_, MU1_EFPGA_TPRAM_COEF_R_ADDR_6_, MU0_EFPGA_TPRAM_OPER_W_DATA_17_, MU0_EFPGA_TPRAM_OPER_W_DATA_16_, MU0_EFPGA_TPRAM_OPER_W_DATA_7_, MU0_EFPGA_TPRAM_OPER_W_DATA_6_, MU0_EFPGA_TPRAM_OPER_W_DATA_15_, MU0_EFPGA_TPRAM_OPER_W_DATA_14_, MU0_EFPGA_TPRAM_OPER_W_DATA_13_, MU0_EFPGA_TPRAM_OPER_W_DATA_12_, MU0_EFPGA_TPRAM_OPER_W_DATA_11_, MU0_EFPGA_TPRAM_OPER_W_DATA_10_, MU0_EFPGA_TPRAM_OPER_W_DATA_9_, MU0_EFPGA_TPRAM_OPER_W_DATA_8_, MU0_EFPGA_TPRAM_OPER_W_DATA_5_, MU0_EFPGA_TPRAM_OPER_W_DATA_4_, MU0_EFPGA_TPRAM_OPER_W_ADDR_8_, MU0_EFPGA_TPRAM_OPER_W_ADDR_7_, MU0_EFPGA_TPRAM_OPER_W_ADDR_6_, MU0_EFPGA_TPRAM_OPER_W_ADDR_5_, MU0_EFPGA_TPRAM_OPER_W_ADDR_4_, MU0_EFPGA_TPRAM_OPER_W_ADDR_3_, MU0_EFPGA_TPRAM_OPER_W_ADDR_2_, MU0_EFPGA_TPRAM_OPER_W_ADDR_1_, MU0_EFPGA_TPRAM_OPER_W_DATA_3_, MU0_EFPGA_TPRAM_OPER_W_DATA_2_, MU0_EFPGA_TPRAM_OPER_W_DATA_1_, MU0_EFPGA_TPRAM_OPER_W_DATA_0_, MU0_EFPGA_TPRAM_OPER_W_CLK, MU0_EFPGA_TPRAM_OPER_W_ADDR_11_, MU0_EFPGA_TPRAM_OPER_W_ADDR_10_, MU0_EFPGA_TPRAM_OPER_W_ADDR_9_, MU0_EFPGA_TPRAM_OPER_W_ADDR_0_, MU0_EFPGA_TPRAM_OPER_WE, MU0_EFPGA_TPRAM_OPER_R_ADDR_7_, MU0_EFPGA_TPRAM_OPER_R_ADDR_6_, MU0_EFPGA_TPRAM_OPER_WDSEL, MU0_EFPGA_TPRAM_OPER_R_MODE_1_, MU0_EFPGA_TPRAM_OPER_R_MODE_0_, MU0_EFPGA_TPRAM_OPER_R_CLK, MU0_EFPGA_TPRAM_OPER_R_ADDR_11_, MU0_EFPGA_TPRAM_OPER_R_ADDR_10_, MU0_EFPGA_TPRAM_OPER_R_ADDR_9_, MU0_EFPGA_TPRAM_OPER_R_ADDR_8_, MU0_EFPGA_TPRAM_OPER_R_ADDR_5_, MU0_EFPGA_TPRAM_OPER_R_ADDR_4_, MU0_EFPGA_MATHB_MAC_OUT_SEL_4_, MU0_EFPGA_MATHB_MAC_OUT_SEL_3_, MU0_EFPGA_MATHB_MAC_OUT_SEL_2_, MU0_EFPGA_MATHB_MAC_OUT_SEL_1_, MU0_EFPGA_MATHB_MAC_OUT_SEL_0_, MU0_EFPGA_MATHB_MAC_ACC_SAT, MU0_EFPGA_MATHB_MAC_ACC_RND, MU0_EFPGA_MATHB_MAC_ACC_CLEAR, MU0_EFPGA_TPRAM_OPER_R_ADDR_3_, MU0_EFPGA_TPRAM_OPER_R_ADDR_2_, MU0_EFPGA_TPRAM_OPER_R_ADDR_1_, MU0_EFPGA_TPRAM_OPER_R_ADDR_0_, MU0_EFPGA_TPRAM_OPER_POWERDN, MU0_EFPGA2MATHB_CLK, MU0_EFPGA_MATHB_CLK_EN, MU0_EFPGA_MATHB_MAC_OUT_SEL_5_, MU0_EFPGA_MATHB_OPER_SEL, MU0_EFPGA_MATHB_OPER_DATA_31_, MU0_EFPGA_MATHB_OPER_DATA_22_, MU0_EFPGA_MATHB_OPER_DATA_21_, MU0_EFPGA_MATHB_OPER_DATA_30_, MU0_EFPGA_MATHB_OPER_DATA_29_, MU0_EFPGA_MATHB_OPER_DATA_28_, MU0_EFPGA_MATHB_OPER_DATA_27_, MU0_EFPGA_MATHB_OPER_DATA_26_, MU0_EFPGA_MATHB_OPER_DATA_25_, MU0_EFPGA_MATHB_OPER_DATA_24_, MU0_EFPGA_MATHB_OPER_DATA_23_, MU0_EFPGA_MATHB_OPER_DATA_20_, MU0_EFPGA_MATHB_OPER_DATA_19_, MU0_EFPGA_MATHB_OPER_DATA_10_, MU0_EFPGA_MATHB_OPER_DATA_9_, MU0_EFPGA_MATHB_OPER_DATA_8_, MU0_EFPGA_MATHB_OPER_DATA_7_, MU0_EFPGA_MATHB_OPER_DATA_6_, MU0_EFPGA_MATHB_OPER_DATA_5_, MU0_EFPGA_MATHB_OPER_DATA_4_, MU0_EFPGA_MATHB_OPER_DATA_3_, MU0_EFPGA_MATHB_OPER_DATA_18_, MU0_EFPGA_MATHB_OPER_DATA_17_, MU0_EFPGA_MATHB_OPER_DATA_16_, MU0_EFPGA_MATHB_OPER_DATA_15_, MU0_EFPGA_MATHB_OPER_DATA_14_, MU0_EFPGA_MATHB_OPER_DATA_13_, MU0_EFPGA_MATHB_OPER_DATA_12_, MU0_EFPGA_MATHB_OPER_DATA_11_, MU0_EFPGA_MATHB_OPER_DATA_2_, MU0_EFPGA_MATHB_OPER_DATA_1_, MU0_EFPGA_MATHB_COEF_DATA_25_, MU0_EFPGA_MATHB_COEF_DATA_24_, MU0_EFPGA_MATHB_OPER_DATA_0_, MU0_EFPGA_MATHB_COEF_SEL, MU0_EFPGA_MATHB_COEF_DATA_31_, MU0_EFPGA_MATHB_COEF_DATA_30_, MU0_EFPGA_MATHB_COEF_DATA_29_, MU0_EFPGA_MATHB_COEF_DATA_28_, MU0_EFPGA_MATHB_COEF_DATA_27_, MU0_EFPGA_MATHB_COEF_DATA_26_, MU1_EFPGA_MATHB_TC_defPin, MU1_EFPGA_MATHB_OPER_defPin_1_, MU1_EFPGA_MATHB_OPER_defPin_0_, MU1_EFPGA_MATHB_COEF_defPin_1_, MU1_EFPGA_MATHB_COEF_defPin_0_, MU0_EFPGA_MATHB_TC_defPin, MU0_EFPGA_MATHB_OPER_defPin_1_, MU0_EFPGA_MATHB_OPER_defPin_0_, MU0_EFPGA_MATHB_COEF_defPin_1_, MU0_EFPGA_MATHB_COEF_defPin_0_, BL_DOUT_0_, BL_DOUT_10_, BL_DOUT_11_, BL_DOUT_12_, BL_DOUT_13_, BL_DOUT_14_, BL_DOUT_15_, BL_DOUT_16_, BL_DOUT_17_, BL_DOUT_18_, BL_DOUT_19_, BL_DOUT_1_, BL_DOUT_20_, BL_DOUT_21_, BL_DOUT_22_, BL_DOUT_23_, BL_DOUT_24_, BL_DOUT_25_, BL_DOUT_26_, BL_DOUT_27_, BL_DOUT_28_, BL_DOUT_29_, BL_DOUT_2_, BL_DOUT_30_, BL_DOUT_31_, BL_DOUT_3_, BL_DOUT_4_, BL_DOUT_5_, BL_DOUT_6_, BL_DOUT_7_, BL_DOUT_8_, BL_DOUT_9_, FB_SPE_OUT_0_, FB_SPE_OUT_1_, FB_SPE_OUT_2_, FB_SPE_OUT_3_, PARALLEL_CFG, supplyBus  );

input   [475:0] supplyBus;

input   CLK0, CLK1, CLK2, CLK3, CLK4, CLK5, fpgaio_data_0_i, fpgaio_data_1_i, fpgaio_data_2_i, fpgaio_data_3_i, fpgaio_data_4_i, fpgaio_data_5_i, fpgaio_data_6_i, fpgaio_data_7_i, udma_cfg_data_8_i, udma_cfg_data_9_i, udma_cfg_data_10_i, udma_cfg_data_11_i, udma_cfg_data_12_i, udma_cfg_data_13_i, udma_cfg_data_14_i, udma_cfg_data_15_i, udma_cfg_data_2_i, udma_cfg_data_3_i, udma_cfg_data_4_i, udma_cfg_data_5_i, udma_cfg_data_6_i, udma_cfg_data_7_i, udma_tx_lin_data_27_i, udma_tx_lin_data_28_i, udma_tx_lin_data_29_i, udma_tx_lin_data_30_i, udma_tx_lin_data_31_i, udma_rx_lin_ready_i, udma_cfg_data_0_i, udma_cfg_data_1_i, udma_tx_lin_data_21_i, udma_tx_lin_data_22_i, udma_tx_lin_data_23_i, udma_tx_lin_data_24_i, udma_tx_lin_data_25_i, udma_tx_lin_data_26_i, udma_tx_lin_data_13_i, udma_tx_lin_data_14_i, udma_tx_lin_data_15_i, udma_tx_lin_data_16_i, udma_tx_lin_data_17_i, udma_tx_lin_data_18_i, udma_tx_lin_data_19_i, udma_tx_lin_data_20_i, udma_tx_lin_data_7_i, udma_tx_lin_data_8_i, udma_tx_lin_data_9_i, udma_tx_lin_data_10_i, udma_tx_lin_data_11_i, udma_tx_lin_data_12_i, udma_tx_lin_valid_i, udma_tx_lin_data_0_i, udma_tx_lin_data_1_i, udma_tx_lin_data_2_i, udma_tx_lin_data_3_i, udma_tx_lin_data_4_i, udma_tx_lin_data_5_i, udma_tx_lin_data_6_i, apb_hwce_pwdata_0_i, apb_hwce_pwdata_1_i, apb_hwce_pwdata_2_i, apb_hwce_pwdata_3_i, apb_hwce_pwdata_4_i, apb_hwce_pwdata_5_i, apb_hwce_pwdata_6_i, apb_hwce_pwdata_7_i, apb_hwce_pwdata_8_i, apb_hwce_pwdata_9_i, apb_hwce_pwdata_10_i, apb_hwce_pwdata_11_i, apb_hwce_pwdata_12_i, apb_hwce_pwdata_13_i, apb_hwce_pwdata_14_i, apb_hwce_pwdata_15_i, apb_hwce_pwdata_16_i, apb_hwce_pwdata_17_i, apb_hwce_pwdata_18_i, apb_hwce_pwdata_19_i, apb_hwce_pwdata_20_i, apb_hwce_pwdata_21_i, apb_hwce_pwdata_22_i, apb_hwce_pwdata_23_i, apb_hwce_pwdata_24_i, apb_hwce_pwdata_25_i, apb_hwce_pwdata_26_i, apb_hwce_pwdata_27_i, apb_hwce_pwdata_28_i, apb_hwce_pwdata_29_i, apb_hwce_pwdata_30_i, apb_hwce_pwdata_31_i, apb_hwce_addr_0_i, apb_hwce_addr_1_i, apb_hwce_addr_2_i, apb_hwce_addr_3_i, apb_hwce_addr_4_i, apb_hwce_addr_5_i, apb_hwce_addr_6_i, apb_hwce_enable_i, apb_hwce_psel_i, apb_hwce_pstrb_i, apb_hwce_pwrite_i, fpgaio_data_28_i, fpgaio_data_29_i, fpgaio_data_30_i, fpgaio_data_31_i, fpgaio_data_32_i, fpgaio_data_33_i, fpgaio_data_34_i, fpgaio_data_35_i, fpgaio_data_36_i, fpgaio_data_37_i, fpgaio_data_38_i, fpgaio_data_39_i, fpgaio_data_40_i, fpgaio_data_41_i, fpgaio_data_42_i, RESET_LB, RESET_LT, fpgaio_data_20_i, fpgaio_data_21_i, fpgaio_data_22_i, fpgaio_data_23_i, fpgaio_data_24_i, fpgaio_data_25_i, fpgaio_data_26_i, fpgaio_data_27_i, udma_cfg_data_30_i, udma_cfg_data_31_i, fpgaio_data_16_i, fpgaio_data_17_i, fpgaio_data_18_i, fpgaio_data_19_i, udma_cfg_data_22_i, udma_cfg_data_23_i, udma_cfg_data_24_i, udma_cfg_data_25_i, udma_cfg_data_26_i, udma_cfg_data_27_i, udma_cfg_data_28_i, udma_cfg_data_29_i, udma_cfg_data_16_i, udma_cfg_data_17_i, udma_cfg_data_18_i, udma_cfg_data_19_i, udma_cfg_data_20_i, udma_cfg_data_21_i, tcdm_r_rdata_p3_8_i, tcdm_r_rdata_p3_9_i, tcdm_r_rdata_p3_10_i, tcdm_r_rdata_p3_11_i, tcdm_r_rdata_p3_12_i, tcdm_r_rdata_p3_13_i, tcdm_r_rdata_p3_14_i, tcdm_r_rdata_p3_15_i, tcdm_r_rdata_p3_2_i, tcdm_r_rdata_p3_3_i, tcdm_r_rdata_p3_4_i, tcdm_r_rdata_p3_5_i, tcdm_r_rdata_p3_6_i, tcdm_r_rdata_p3_7_i, tcdm_r_rdata_p2_28_i, tcdm_r_rdata_p2_29_i, tcdm_r_rdata_p2_30_i, tcdm_r_rdata_p2_31_i, tcdm_gnt_p2_i, tcdm_r_valid_p2_i, tcdm_r_rdata_p3_0_i, tcdm_r_rdata_p3_1_i, tcdm_r_rdata_p2_22_i, tcdm_r_rdata_p2_23_i, tcdm_r_rdata_p2_24_i, tcdm_r_rdata_p2_25_i, tcdm_r_rdata_p2_26_i, tcdm_r_rdata_p2_27_i, tcdm_r_rdata_p2_14_i, tcdm_r_rdata_p2_15_i, tcdm_r_rdata_p2_16_i, tcdm_r_rdata_p2_17_i, tcdm_r_rdata_p2_18_i, tcdm_r_rdata_p2_19_i, tcdm_r_rdata_p2_20_i, tcdm_r_rdata_p2_21_i, tcdm_r_rdata_p2_8_i, tcdm_r_rdata_p2_9_i, tcdm_r_rdata_p2_10_i, tcdm_r_rdata_p2_11_i, tcdm_r_rdata_p2_12_i, tcdm_r_rdata_p2_13_i, tcdm_r_rdata_p2_0_i, tcdm_r_rdata_p2_1_i, tcdm_r_rdata_p2_2_i, tcdm_r_rdata_p2_3_i, tcdm_r_rdata_p2_4_i, tcdm_r_rdata_p2_5_i, tcdm_r_rdata_p2_6_i, tcdm_r_rdata_p2_7_i, tcdm_r_rdata_p0_0_i, tcdm_r_rdata_p0_1_i, tcdm_r_rdata_p0_2_i, tcdm_r_rdata_p0_3_i, tcdm_r_rdata_p0_4_i, tcdm_r_rdata_p0_5_i, tcdm_r_rdata_p0_6_i, tcdm_r_rdata_p0_7_i, tcdm_r_rdata_p0_8_i, tcdm_r_rdata_p0_9_i, tcdm_r_rdata_p0_10_i, tcdm_r_rdata_p0_11_i, tcdm_r_rdata_p0_12_i, tcdm_r_rdata_p0_13_i, tcdm_r_rdata_p0_14_i, tcdm_r_rdata_p0_15_i, tcdm_r_rdata_p0_16_i, tcdm_r_rdata_p0_17_i, tcdm_r_rdata_p0_18_i, tcdm_r_rdata_p0_19_i, tcdm_r_rdata_p0_20_i, tcdm_r_rdata_p0_21_i, tcdm_r_rdata_p0_22_i, tcdm_r_rdata_p0_23_i, tcdm_r_rdata_p0_24_i, tcdm_r_rdata_p0_25_i, tcdm_r_rdata_p0_26_i, tcdm_r_rdata_p0_27_i, tcdm_r_rdata_p0_28_i, tcdm_r_rdata_p0_29_i, tcdm_r_rdata_p0_30_i, tcdm_r_rdata_p0_31_i, tcdm_gnt_p0_i, tcdm_r_valid_p0_i, tcdm_r_rdata_p1_0_i, tcdm_r_rdata_p1_1_i, tcdm_r_rdata_p1_2_i, tcdm_r_rdata_p1_3_i, tcdm_r_rdata_p1_4_i, tcdm_r_rdata_p1_5_i, tcdm_r_rdata_p1_6_i, tcdm_r_rdata_p1_7_i, tcdm_r_rdata_p1_8_i, tcdm_r_rdata_p1_9_i, tcdm_r_rdata_p1_10_i, tcdm_r_rdata_p1_11_i, tcdm_r_rdata_p1_12_i, tcdm_r_rdata_p1_13_i, tcdm_r_rdata_p1_14_i, tcdm_r_rdata_p1_15_i, tcdm_r_rdata_p1_16_i, tcdm_r_rdata_p1_17_i, tcdm_r_rdata_p1_18_i, tcdm_r_rdata_p1_19_i, tcdm_r_rdata_p1_20_i, tcdm_r_rdata_p1_21_i, tcdm_r_rdata_p1_22_i, tcdm_r_rdata_p1_23_i, tcdm_r_rdata_p1_24_i, tcdm_r_rdata_p1_25_i, tcdm_r_rdata_p1_26_i, tcdm_r_rdata_p1_27_i, tcdm_r_rdata_p1_28_i, tcdm_r_rdata_p1_29_i, tcdm_r_rdata_p1_30_i, tcdm_r_rdata_p1_31_i, tcdm_gnt_p1_i, tcdm_r_valid_p1_i, fpgaio_data_8_i, fpgaio_data_9_i, fpgaio_data_10_i, fpgaio_data_11_i, RESET_RB, fpgaio_data_14_i, fpgaio_data_15_i, RESET_RT, tcdm_r_rdata_p3_30_i, tcdm_r_rdata_p3_31_i, tcdm_gnt_p3_i, tcdm_r_valid_p3_i, fpgaio_data_12_i, fpgaio_data_13_i, tcdm_r_rdata_p3_22_i, tcdm_r_rdata_p3_23_i, tcdm_r_rdata_p3_24_i, tcdm_r_rdata_p3_25_i, tcdm_r_rdata_p3_26_i, tcdm_r_rdata_p3_27_i, tcdm_r_rdata_p3_28_i, tcdm_r_rdata_p3_29_i, tcdm_r_rdata_p3_16_i, tcdm_r_rdata_p3_17_i, tcdm_r_rdata_p3_18_i, tcdm_r_rdata_p3_19_i, tcdm_r_rdata_p3_20_i, tcdm_r_rdata_p3_21_i, MU0_MATHB_EFPGA_MAC_OUT_7_, MU0_MATHB_EFPGA_MAC_OUT_6_, MU0_MATHB_EFPGA_MAC_OUT_5_, MU0_MATHB_EFPGA_MAC_OUT_4_, MU0_MATHB_EFPGA_MAC_OUT_3_, MU0_MATHB_EFPGA_MAC_OUT_2_, MU0_MATHB_EFPGA_MAC_OUT_1_, MU0_MATHB_EFPGA_MAC_OUT_0_, MU0_TPRAM_EFPGA_COEF_R_DATA_31_, MU0_TPRAM_EFPGA_COEF_R_DATA_30_, MU0_TPRAM_EFPGA_COEF_R_DATA_29_, MU0_TPRAM_EFPGA_COEF_R_DATA_28_, MU0_TPRAM_EFPGA_COEF_R_DATA_27_, MU0_TPRAM_EFPGA_COEF_R_DATA_26_, MU0_TPRAM_EFPGA_COEF_R_DATA_25_, MU0_TPRAM_EFPGA_COEF_R_DATA_24_, MU0_TPRAM_EFPGA_COEF_R_DATA_23_, MU0_TPRAM_EFPGA_COEF_R_DATA_22_, MU0_TPRAM_EFPGA_COEF_R_DATA_21_, MU0_TPRAM_EFPGA_COEF_R_DATA_20_, MU0_TPRAM_EFPGA_COEF_R_DATA_19_, MU0_TPRAM_EFPGA_COEF_R_DATA_18_, MU0_TPRAM_EFPGA_COEF_R_DATA_17_, MU0_TPRAM_EFPGA_COEF_R_DATA_16_, MU0_TPRAM_EFPGA_COEF_R_DATA_15_, MU0_TPRAM_EFPGA_COEF_R_DATA_14_, MU0_TPRAM_EFPGA_COEF_R_DATA_13_, MU0_TPRAM_EFPGA_COEF_R_DATA_12_, MU0_TPRAM_EFPGA_COEF_R_DATA_11_, MU0_TPRAM_EFPGA_COEF_R_DATA_10_, MU0_TPRAM_EFPGA_COEF_R_DATA_9_, MU0_TPRAM_EFPGA_COEF_R_DATA_8_, MU0_TPRAM_EFPGA_COEF_R_DATA_7_, MU0_TPRAM_EFPGA_COEF_R_DATA_6_, MU0_TPRAM_EFPGA_COEF_R_DATA_5_, MU0_TPRAM_EFPGA_COEF_R_DATA_4_, MU0_TPRAM_EFPGA_COEF_R_DATA_3_, MU0_TPRAM_EFPGA_COEF_R_DATA_2_, MU0_TPRAM_EFPGA_COEF_R_DATA_1_, MU0_TPRAM_EFPGA_COEF_R_DATA_0_, MU1_TPRAM_EFPGA_OPER_R_DATA_31_, MU1_TPRAM_EFPGA_OPER_R_DATA_30_, MU1_TPRAM_EFPGA_OPER_R_DATA_29_, MU1_TPRAM_EFPGA_OPER_R_DATA_28_, MU1_TPRAM_EFPGA_OPER_R_DATA_27_, MU1_TPRAM_EFPGA_OPER_R_DATA_26_, MU1_TPRAM_EFPGA_OPER_R_DATA_25_, MU1_TPRAM_EFPGA_OPER_R_DATA_24_, MU1_TPRAM_EFPGA_OPER_R_DATA_23_, MU1_TPRAM_EFPGA_OPER_R_DATA_22_, MU1_TPRAM_EFPGA_OPER_R_DATA_21_, MU1_TPRAM_EFPGA_OPER_R_DATA_20_, MU1_TPRAM_EFPGA_OPER_R_DATA_19_, MU1_TPRAM_EFPGA_OPER_R_DATA_18_, MU1_TPRAM_EFPGA_OPER_R_DATA_17_, MU1_TPRAM_EFPGA_OPER_R_DATA_16_, MU1_TPRAM_EFPGA_OPER_R_DATA_15_, MU1_TPRAM_EFPGA_OPER_R_DATA_14_, MU1_TPRAM_EFPGA_OPER_R_DATA_13_, MU1_TPRAM_EFPGA_OPER_R_DATA_12_, MU0_TPRAM_EFPGA_OPER_R_DATA_31_, MU0_TPRAM_EFPGA_OPER_R_DATA_30_, MU0_TPRAM_EFPGA_OPER_R_DATA_29_, MU0_TPRAM_EFPGA_OPER_R_DATA_28_, MU1_TPRAM_EFPGA_OPER_R_DATA_11_, MU1_TPRAM_EFPGA_OPER_R_DATA_10_, MU1_TPRAM_EFPGA_OPER_R_DATA_9_, MU1_TPRAM_EFPGA_OPER_R_DATA_8_, MU1_TPRAM_EFPGA_OPER_R_DATA_7_, MU1_TPRAM_EFPGA_OPER_R_DATA_6_, MU1_TPRAM_EFPGA_OPER_R_DATA_5_, MU1_TPRAM_EFPGA_OPER_R_DATA_4_, MU1_TPRAM_EFPGA_OPER_R_DATA_3_, MU1_TPRAM_EFPGA_OPER_R_DATA_2_, MU1_TPRAM_EFPGA_OPER_R_DATA_1_, MU1_TPRAM_EFPGA_OPER_R_DATA_0_, MU1_MATHB_EFPGA_MAC_OUT_31_, MU1_MATHB_EFPGA_MAC_OUT_30_, MU1_MATHB_EFPGA_MAC_OUT_29_, MU1_MATHB_EFPGA_MAC_OUT_28_, MU1_MATHB_EFPGA_MAC_OUT_27_, MU1_MATHB_EFPGA_MAC_OUT_26_, MU1_MATHB_EFPGA_MAC_OUT_25_, MU1_MATHB_EFPGA_MAC_OUT_24_, MU1_MATHB_EFPGA_MAC_OUT_23_, MU1_MATHB_EFPGA_MAC_OUT_22_, MU1_MATHB_EFPGA_MAC_OUT_21_, MU1_MATHB_EFPGA_MAC_OUT_20_, MU1_MATHB_EFPGA_MAC_OUT_19_, MU1_MATHB_EFPGA_MAC_OUT_18_, MU1_MATHB_EFPGA_MAC_OUT_17_, MU1_MATHB_EFPGA_MAC_OUT_16_, MU1_MATHB_EFPGA_MAC_OUT_15_, MU1_MATHB_EFPGA_MAC_OUT_14_, MU1_MATHB_EFPGA_MAC_OUT_13_, MU1_MATHB_EFPGA_MAC_OUT_12_, MU1_MATHB_EFPGA_MAC_OUT_11_, MU1_MATHB_EFPGA_MAC_OUT_10_, MU1_MATHB_EFPGA_MAC_OUT_9_, MU1_MATHB_EFPGA_MAC_OUT_8_, MU1_MATHB_EFPGA_MAC_OUT_7_, MU1_MATHB_EFPGA_MAC_OUT_6_, MU1_MATHB_EFPGA_MAC_OUT_5_, MU1_MATHB_EFPGA_MAC_OUT_4_, MU1_MATHB_EFPGA_MAC_OUT_3_, MU1_MATHB_EFPGA_MAC_OUT_2_, MU1_MATHB_EFPGA_MAC_OUT_1_, MU1_MATHB_EFPGA_MAC_OUT_0_, MU1_TPRAM_EFPGA_COEF_R_DATA_31_, MU1_TPRAM_EFPGA_COEF_R_DATA_30_, MU1_TPRAM_EFPGA_COEF_R_DATA_29_, MU1_TPRAM_EFPGA_COEF_R_DATA_28_, MU1_TPRAM_EFPGA_COEF_R_DATA_27_, MU1_TPRAM_EFPGA_COEF_R_DATA_26_, MU1_TPRAM_EFPGA_COEF_R_DATA_25_, MU1_TPRAM_EFPGA_COEF_R_DATA_24_, MU1_TPRAM_EFPGA_COEF_R_DATA_23_, MU1_TPRAM_EFPGA_COEF_R_DATA_22_, MU1_TPRAM_EFPGA_COEF_R_DATA_21_, MU1_TPRAM_EFPGA_COEF_R_DATA_20_, MU1_TPRAM_EFPGA_COEF_R_DATA_19_, MU1_TPRAM_EFPGA_COEF_R_DATA_18_, MU0_TPRAM_EFPGA_OPER_R_DATA_27_, MU0_TPRAM_EFPGA_OPER_R_DATA_26_, MU0_TPRAM_EFPGA_OPER_R_DATA_25_, MU0_TPRAM_EFPGA_OPER_R_DATA_24_, MU0_TPRAM_EFPGA_OPER_R_DATA_23_, MU0_TPRAM_EFPGA_OPER_R_DATA_22_, MU0_TPRAM_EFPGA_OPER_R_DATA_21_, MU0_TPRAM_EFPGA_OPER_R_DATA_20_, MU1_TPRAM_EFPGA_COEF_R_DATA_17_, MU1_TPRAM_EFPGA_COEF_R_DATA_16_, MU1_TPRAM_EFPGA_COEF_R_DATA_15_, MU1_TPRAM_EFPGA_COEF_R_DATA_14_, MU1_TPRAM_EFPGA_COEF_R_DATA_13_, MU1_TPRAM_EFPGA_COEF_R_DATA_12_, MU1_TPRAM_EFPGA_COEF_R_DATA_11_, MU1_TPRAM_EFPGA_COEF_R_DATA_10_, MU1_TPRAM_EFPGA_COEF_R_DATA_9_, MU1_TPRAM_EFPGA_COEF_R_DATA_8_, MU1_TPRAM_EFPGA_COEF_R_DATA_7_, MU1_TPRAM_EFPGA_COEF_R_DATA_6_, MU1_TPRAM_EFPGA_COEF_R_DATA_5_, MU1_TPRAM_EFPGA_COEF_R_DATA_4_, MU1_TPRAM_EFPGA_COEF_R_DATA_3_, MU1_TPRAM_EFPGA_COEF_R_DATA_2_, MU1_TPRAM_EFPGA_COEF_R_DATA_1_, MU1_TPRAM_EFPGA_COEF_R_DATA_0_, MU0_TPRAM_EFPGA_OPER_R_DATA_19_, MU0_TPRAM_EFPGA_OPER_R_DATA_18_, MU0_TPRAM_EFPGA_OPER_R_DATA_17_, MU0_TPRAM_EFPGA_OPER_R_DATA_16_, MU0_TPRAM_EFPGA_OPER_R_DATA_15_, MU0_TPRAM_EFPGA_OPER_R_DATA_14_, MU0_TPRAM_EFPGA_OPER_R_DATA_13_, MU0_TPRAM_EFPGA_OPER_R_DATA_12_, MU0_TPRAM_EFPGA_OPER_R_DATA_11_, MU0_TPRAM_EFPGA_OPER_R_DATA_10_, MU0_TPRAM_EFPGA_OPER_R_DATA_9_, MU0_TPRAM_EFPGA_OPER_R_DATA_8_, MU0_TPRAM_EFPGA_OPER_R_DATA_7_, MU0_TPRAM_EFPGA_OPER_R_DATA_6_, MU0_TPRAM_EFPGA_OPER_R_DATA_5_, MU0_TPRAM_EFPGA_OPER_R_DATA_4_, MU0_TPRAM_EFPGA_OPER_R_DATA_3_, MU0_TPRAM_EFPGA_OPER_R_DATA_2_, MU0_TPRAM_EFPGA_OPER_R_DATA_1_, MU0_TPRAM_EFPGA_OPER_R_DATA_0_, MU0_MATHB_EFPGA_MAC_OUT_31_, MU0_MATHB_EFPGA_MAC_OUT_30_, MU0_MATHB_EFPGA_MAC_OUT_29_, MU0_MATHB_EFPGA_MAC_OUT_28_, MU0_MATHB_EFPGA_MAC_OUT_27_, MU0_MATHB_EFPGA_MAC_OUT_26_, MU0_MATHB_EFPGA_MAC_OUT_25_, MU0_MATHB_EFPGA_MAC_OUT_24_, MU0_MATHB_EFPGA_MAC_OUT_23_, MU0_MATHB_EFPGA_MAC_OUT_22_, MU0_MATHB_EFPGA_MAC_OUT_21_, MU0_MATHB_EFPGA_MAC_OUT_20_, MU0_MATHB_EFPGA_MAC_OUT_19_, MU0_MATHB_EFPGA_MAC_OUT_18_, MU0_MATHB_EFPGA_MAC_OUT_17_, MU0_MATHB_EFPGA_MAC_OUT_16_, MU0_MATHB_EFPGA_MAC_OUT_15_, MU0_MATHB_EFPGA_MAC_OUT_14_, MU0_MATHB_EFPGA_MAC_OUT_13_, MU0_MATHB_EFPGA_MAC_OUT_12_, MU0_MATHB_EFPGA_MAC_OUT_11_, MU0_MATHB_EFPGA_MAC_OUT_10_, MU0_MATHB_EFPGA_MAC_OUT_9_, MU0_MATHB_EFPGA_MAC_OUT_8_,  M_0_, BL_CLK, BL_DIN_0_, BL_DIN_10_, BL_DIN_11_, BL_DIN_12_, BL_DIN_13_, BL_DIN_14_, BL_DIN_15_, BL_DIN_16_, BL_DIN_17_, BL_DIN_18_, BL_DIN_19_, BL_DIN_1_, BL_DIN_20_, BL_DIN_21_, BL_DIN_22_, BL_DIN_23_, BL_DIN_24_, BL_DIN_25_, BL_DIN_26_, BL_DIN_27_, BL_DIN_28_, BL_DIN_29_, BL_DIN_2_, BL_DIN_30_, BL_DIN_31_, BL_DIN_3_, BL_DIN_4_, BL_DIN_5_, BL_DIN_6_, BL_DIN_7_, BL_DIN_8_, BL_DIN_9_, BL_PWRGATE_0_, BL_PWRGATE_1_, BL_PWRGATE_2_, BL_PWRGATE_3_, CLOAD_DIN_SEL, DIN_INT_L_ONLY, DIN_INT_R_ONLY, DIN_SLC_TB_INT, FB_CFG_DONE, FB_ISO_ENB, FB_SPE_IN_0_, FB_SPE_IN_1_, FB_SPE_IN_2_, FB_SPE_IN_3_, ISO_EN_0_, ISO_EN_1_, ISO_EN_2_, ISO_EN_3_, MLATCH, M_1_, M_2_, M_3_, M_4_, M_5_, NB, PB, PCHG_B, PI_PWR_0_, PI_PWR_1_, PI_PWR_2_, PI_PWR_3_, POR, PROG_0_, PROG_1_, PROG_2_, PROG_3_, PROG_IFX, PWR_GATE, RE, STM, VLP_CLKDIS_0_, VLP_CLKDIS_1_, VLP_CLKDIS_2_, VLP_CLKDIS_3_, VLP_CLKDIS_IFX, VLP_PWRDIS_0_, VLP_PWRDIS_1_, VLP_PWRDIS_2_, VLP_PWRDIS_3_, VLP_PWRDIS_IFX, VLP_SRDIS_0_, VLP_SRDIS_1_, VLP_SRDIS_2_, VLP_SRDIS_3_, VLP_SRDIS_IFX, WE, WE_INT, WL_CLK, WL_CLOAD_SEL_0_, WL_CLOAD_SEL_1_, WL_CLOAD_SEL_2_, WL_DIN_0_, WL_DIN_1_, WL_DIN_2_, WL_DIN_3_, WL_DIN_4_, WL_DIN_5_, WL_EN, WL_INT_DIN_SEL, WL_PWRGATE_0_, WL_PWRGATE_1_, WL_RESETB, WL_SEL_0_, WL_SEL_1_, WL_SEL_2_, WL_SEL_3_, WL_SEL_TB_INT;


output   fpgaio_oe_0_o, fpgaio_data_0_o, fpgaio_oe_1_o, fpgaio_data_1_o, fpgaio_oe_2_o, fpgaio_data_2_o, fpgaio_oe_3_o, fpgaio_data_3_o, fpgaio_oe_4_o, fpgaio_data_4_o, fpgaio_oe_5_o, fpgaio_data_5_o, fpgaio_oe_6_o, fpgaio_data_6_o, fpgaio_oe_7_o, fpgaio_data_7_o, fpgaio_oe_20_o, fpgaio_data_20_o, fpgaio_oe_25_o, fpgaio_data_25_o, fpgaio_oe_26_o, fpgaio_data_26_o, fpgaio_oe_27_o, fpgaio_data_27_o, fpgaio_oe_21_o, fpgaio_data_21_o, fpgaio_oe_22_o, fpgaio_data_22_o, fpgaio_oe_23_o, fpgaio_data_23_o, fpgaio_oe_24_o, fpgaio_data_24_o, events_12_o, events_13_o, fpgaio_oe_19_o, fpgaio_data_19_o, events_14_o, events_15_o, fpgaio_oe_16_o, fpgaio_data_16_o, fpgaio_oe_17_o, fpgaio_data_17_o, fpgaio_oe_18_o, fpgaio_data_18_o, udma_cfg_data_26_o, udma_cfg_data_27_o, events_4_o, events_5_o, events_6_o, events_7_o, events_8_o, events_9_o, events_10_o, events_11_o, udma_cfg_data_28_o, udma_cfg_data_29_o, udma_cfg_data_30_o, udma_cfg_data_31_o, events_0_o, events_1_o, events_2_o, events_3_o, udma_cfg_data_14_o, udma_cfg_data_15_o, udma_cfg_data_24_o, udma_cfg_data_25_o, udma_cfg_data_16_o, udma_cfg_data_17_o, udma_cfg_data_18_o, udma_cfg_data_19_o, udma_cfg_data_20_o, udma_cfg_data_21_o, udma_cfg_data_22_o, udma_cfg_data_23_o, udma_rx_lin_data_28_o, udma_rx_lin_data_29_o, udma_cfg_data_6_o, udma_cfg_data_7_o, udma_cfg_data_8_o, udma_cfg_data_9_o, udma_cfg_data_10_o, udma_cfg_data_11_o, udma_cfg_data_12_o, udma_cfg_data_13_o, udma_rx_lin_data_30_o, udma_rx_lin_data_31_o, udma_cfg_data_0_o, udma_cfg_data_1_o, udma_cfg_data_2_o, udma_cfg_data_3_o, udma_cfg_data_4_o, udma_cfg_data_5_o, udma_rx_lin_data_16_o, udma_rx_lin_data_17_o, udma_rx_lin_data_26_o, udma_rx_lin_data_27_o, udma_rx_lin_data_18_o, udma_rx_lin_data_19_o, udma_rx_lin_data_20_o, udma_rx_lin_data_21_o, udma_rx_lin_data_22_o, udma_rx_lin_data_23_o, udma_rx_lin_data_24_o, udma_rx_lin_data_25_o, udma_tx_lin_ready_o, udma_rx_lin_valid_o, udma_rx_lin_data_8_o, udma_rx_lin_data_9_o, udma_rx_lin_data_10_o, udma_rx_lin_data_11_o, udma_rx_lin_data_12_o, udma_rx_lin_data_13_o, udma_rx_lin_data_14_o, udma_rx_lin_data_15_o, udma_rx_lin_data_0_o, udma_rx_lin_data_1_o, udma_rx_lin_data_2_o, udma_rx_lin_data_3_o, udma_rx_lin_data_4_o, udma_rx_lin_data_5_o, udma_rx_lin_data_6_o, udma_rx_lin_data_7_o, apb_hwce_prdata_0_o, apb_hwce_prdata_1_o, apb_hwce_prdata_10_o, apb_hwce_prdata_11_o, apb_hwce_prdata_2_o, apb_hwce_prdata_3_o, apb_hwce_prdata_4_o, apb_hwce_prdata_5_o, apb_hwce_prdata_6_o, apb_hwce_prdata_7_o, apb_hwce_prdata_8_o, apb_hwce_prdata_9_o, apb_hwce_prdata_12_o, apb_hwce_prdata_13_o, apb_hwce_prdata_22_o, apb_hwce_prdata_23_o, apb_hwce_prdata_24_o, apb_hwce_prdata_25_o, apb_hwce_prdata_26_o, apb_hwce_prdata_27_o, apb_hwce_prdata_28_o, apb_hwce_prdata_29_o, apb_hwce_prdata_14_o, apb_hwce_prdata_15_o, apb_hwce_prdata_16_o, apb_hwce_prdata_17_o, apb_hwce_prdata_18_o, apb_hwce_prdata_19_o, apb_hwce_prdata_20_o, apb_hwce_prdata_21_o, apb_hwce_prdata_30_o, apb_hwce_prdata_31_o, fpgaio_oe_31_o, fpgaio_data_31_o, apb_hwce_ready_o, apb_hwce_pslverr_o, fpgaio_oe_28_o, fpgaio_data_28_o, fpgaio_oe_29_o, fpgaio_data_29_o, fpgaio_oe_30_o, fpgaio_data_30_o, fpgaio_oe_32_o, fpgaio_data_32_o, fpgaio_oe_37_o, fpgaio_data_37_o, fpgaio_oe_38_o, fpgaio_data_38_o, fpgaio_oe_39_o, fpgaio_data_39_o, fpgaio_oe_40_o, fpgaio_data_40_o, fpgaio_oe_33_o, fpgaio_data_33_o, fpgaio_oe_34_o, fpgaio_data_34_o, fpgaio_oe_35_o, fpgaio_data_35_o, fpgaio_oe_36_o, fpgaio_data_36_o, fpgaio_oe_41_o, fpgaio_data_41_o, fpgaio_oe_42_o, fpgaio_data_42_o, tcdm_addr_p3_16_o, tcdm_wdata_p3_16_o, tcdm_wdata_p3_22_o, tcdm_wdata_p3_23_o, tcdm_wdata_p3_24_o, tcdm_wdata_p3_25_o, tcdm_wdata_p3_26_o, tcdm_wdata_p3_27_o, tcdm_wdata_p3_28_o, tcdm_wdata_p3_29_o, tcdm_addr_p3_17_o, tcdm_wdata_p3_17_o, tcdm_addr_p3_18_o, tcdm_wdata_p3_18_o, tcdm_addr_p3_19_o, tcdm_wdata_p3_19_o, tcdm_wdata_p3_20_o, tcdm_wdata_p3_21_o, tcdm_addr_p3_10_o, tcdm_wdata_p3_10_o, tcdm_addr_p3_15_o, tcdm_wdata_p3_15_o, tcdm_addr_p3_11_o, tcdm_wdata_p3_11_o, tcdm_addr_p3_12_o, tcdm_wdata_p3_12_o, tcdm_addr_p3_13_o, tcdm_wdata_p3_13_o, tcdm_addr_p3_14_o, tcdm_wdata_p3_14_o, tcdm_addr_p3_1_o, tcdm_wdata_p3_1_o, tcdm_addr_p3_6_o, tcdm_wdata_p3_6_o, tcdm_addr_p3_7_o, tcdm_wdata_p3_7_o, tcdm_addr_p3_8_o, tcdm_wdata_p3_8_o, tcdm_addr_p3_9_o, tcdm_wdata_p3_9_o, tcdm_addr_p3_2_o, tcdm_wdata_p3_2_o, tcdm_addr_p3_3_o, tcdm_wdata_p3_3_o, tcdm_addr_p3_4_o, tcdm_wdata_p3_4_o, tcdm_addr_p3_5_o, tcdm_wdata_p3_5_o, tcdm_wdata_p2_28_o, tcdm_wdata_p2_29_o, tcdm_addr_p3_0_o, tcdm_wdata_p3_0_o, tcdm_wdata_p2_30_o, tcdm_wdata_p2_31_o, tcdm_req_p2_o, tcdm_wen_p2_o, tcdm_be_p2_0_o, tcdm_be_p2_1_o, tcdm_be_p2_2_o, tcdm_be_p2_3_o, tcdm_addr_p2_15_o, tcdm_wdata_p2_15_o, tcdm_wdata_p2_20_o, tcdm_wdata_p2_21_o, tcdm_wdata_p2_22_o, tcdm_wdata_p2_23_o, tcdm_wdata_p2_24_o, tcdm_wdata_p2_25_o, tcdm_wdata_p2_26_o, tcdm_wdata_p2_27_o, tcdm_addr_p2_16_o, tcdm_wdata_p2_16_o, tcdm_addr_p2_17_o, tcdm_wdata_p2_17_o, tcdm_addr_p2_18_o, tcdm_wdata_p2_18_o, tcdm_addr_p2_19_o, tcdm_wdata_p2_19_o, tcdm_addr_p2_9_o, tcdm_wdata_p2_9_o, tcdm_addr_p2_14_o, tcdm_wdata_p2_14_o, tcdm_addr_p2_10_o, tcdm_wdata_p2_10_o, tcdm_addr_p2_11_o, tcdm_wdata_p2_11_o, tcdm_addr_p2_12_o, tcdm_wdata_p2_12_o, tcdm_addr_p2_13_o, tcdm_wdata_p2_13_o, tcdm_addr_p2_0_o, tcdm_wdata_p2_0_o, tcdm_addr_p2_5_o, tcdm_wdata_p2_5_o, tcdm_addr_p2_6_o, tcdm_wdata_p2_6_o, tcdm_addr_p2_7_o, tcdm_wdata_p2_7_o, tcdm_addr_p2_8_o, tcdm_wdata_p2_8_o, tcdm_addr_p2_1_o, tcdm_wdata_p2_1_o, tcdm_addr_p2_2_o, tcdm_wdata_p2_2_o, tcdm_addr_p2_3_o, tcdm_wdata_p2_3_o, tcdm_addr_p2_4_o, tcdm_wdata_p2_4_o, tcdm_addr_p0_0_o, tcdm_wdata_p0_0_o, tcdm_addr_p0_5_o, tcdm_wdata_p0_5_o, tcdm_addr_p0_1_o, tcdm_wdata_p0_1_o, tcdm_addr_p0_2_o, tcdm_wdata_p0_2_o, tcdm_addr_p0_3_o, tcdm_wdata_p0_3_o, tcdm_addr_p0_4_o, tcdm_wdata_p0_4_o, tcdm_addr_p0_6_o, tcdm_wdata_p0_6_o, tcdm_addr_p0_11_o, tcdm_wdata_p0_11_o, tcdm_addr_p0_12_o, tcdm_wdata_p0_12_o, tcdm_addr_p0_13_o, tcdm_wdata_p0_13_o, tcdm_addr_p0_14_o, tcdm_wdata_p0_14_o, tcdm_addr_p0_7_o, tcdm_wdata_p0_7_o, tcdm_addr_p0_8_o, tcdm_wdata_p0_8_o, tcdm_addr_p0_9_o, tcdm_wdata_p0_9_o, tcdm_addr_p0_10_o, tcdm_wdata_p0_10_o, tcdm_addr_p0_15_o, tcdm_wdata_p0_15_o, tcdm_wdata_p0_20_o, tcdm_wdata_p0_21_o, tcdm_addr_p0_16_o, tcdm_wdata_p0_16_o, tcdm_addr_p0_17_o, tcdm_wdata_p0_17_o, tcdm_addr_p0_18_o, tcdm_wdata_p0_18_o, tcdm_addr_p0_19_o, tcdm_wdata_p0_19_o, tcdm_wdata_p0_22_o, tcdm_wdata_p0_23_o, tcdm_req_p0_o, tcdm_wen_p0_o, tcdm_be_p0_0_o, tcdm_be_p0_1_o, tcdm_be_p0_2_o, tcdm_be_p0_3_o, tcdm_addr_p1_0_o, tcdm_wdata_p1_0_o, tcdm_wdata_p0_24_o, tcdm_wdata_p0_25_o, tcdm_wdata_p0_26_o, tcdm_wdata_p0_27_o, tcdm_wdata_p0_28_o, tcdm_wdata_p0_29_o, tcdm_wdata_p0_30_o, tcdm_wdata_p0_31_o, tcdm_addr_p1_1_o, tcdm_wdata_p1_1_o, tcdm_addr_p1_6_o, tcdm_wdata_p1_6_o, tcdm_addr_p1_2_o, tcdm_wdata_p1_2_o, tcdm_addr_p1_3_o, tcdm_wdata_p1_3_o, tcdm_addr_p1_4_o, tcdm_wdata_p1_4_o, tcdm_addr_p1_5_o, tcdm_wdata_p1_5_o, tcdm_addr_p1_7_o, tcdm_wdata_p1_7_o, tcdm_addr_p1_12_o, tcdm_wdata_p1_12_o, tcdm_addr_p1_13_o, tcdm_wdata_p1_13_o, tcdm_addr_p1_14_o, tcdm_wdata_p1_14_o, tcdm_addr_p1_15_o, tcdm_wdata_p1_15_o, tcdm_addr_p1_8_o, tcdm_wdata_p1_8_o, tcdm_addr_p1_9_o, tcdm_wdata_p1_9_o, tcdm_addr_p1_10_o, tcdm_wdata_p1_10_o, tcdm_addr_p1_11_o, tcdm_wdata_p1_11_o, tcdm_addr_p1_16_o, tcdm_wdata_p1_16_o, tcdm_wdata_p1_22_o, tcdm_wdata_p1_23_o, tcdm_addr_p1_17_o, tcdm_wdata_p1_17_o, tcdm_addr_p1_18_o, tcdm_wdata_p1_18_o, tcdm_addr_p1_19_o, tcdm_wdata_p1_19_o, tcdm_wdata_p1_20_o, tcdm_wdata_p1_21_o, tcdm_wdata_p1_24_o, tcdm_wdata_p1_25_o, tcdm_be_p1_0_o, tcdm_be_p1_1_o, tcdm_be_p1_2_o, tcdm_be_p1_3_o, fpgaio_oe_8_o, fpgaio_data_8_o, fpgaio_oe_9_o, fpgaio_data_9_o, tcdm_wdata_p1_26_o, tcdm_wdata_p1_27_o, tcdm_wdata_p1_28_o, tcdm_wdata_p1_29_o, tcdm_wdata_p1_30_o, tcdm_wdata_p1_31_o, tcdm_req_p1_o, tcdm_wen_p1_o, fpgaio_oe_10_o, fpgaio_data_10_o, fpgaio_oe_11_o, fpgaio_data_11_o, fpgaio_oe_14_o, fpgaio_data_14_o, fpgaio_oe_15_o, fpgaio_data_15_o, tcdm_wdata_p3_30_o, tcdm_wdata_p3_31_o, fpgaio_oe_13_o, fpgaio_data_13_o, tcdm_req_p3_o, tcdm_wen_p3_o, tcdm_be_p3_0_o, tcdm_be_p3_1_o, tcdm_be_p3_2_o, tcdm_be_p3_3_o, fpgaio_oe_12_o, fpgaio_data_12_o, MU0_EFPGA_MATHB_COEF_DATA_23_, MU0_EFPGA_MATHB_COEF_DATA_22_, MU0_EFPGA_MATHB_COEF_DATA_13_, MU0_EFPGA_MATHB_COEF_DATA_12_, MU0_EFPGA_MATHB_COEF_DATA_11_, MU0_EFPGA_MATHB_COEF_DATA_10_, MU0_EFPGA_MATHB_COEF_DATA_9_, MU0_EFPGA_MATHB_COEF_DATA_8_, MU0_EFPGA_MATHB_COEF_DATA_7_, MU0_EFPGA_MATHB_COEF_DATA_6_, MU0_EFPGA_MATHB_COEF_DATA_21_, MU0_EFPGA_MATHB_COEF_DATA_20_, MU0_EFPGA_MATHB_COEF_DATA_19_, MU0_EFPGA_MATHB_COEF_DATA_18_, MU0_EFPGA_MATHB_COEF_DATA_17_, MU0_EFPGA_MATHB_COEF_DATA_16_, MU0_EFPGA_MATHB_COEF_DATA_15_, MU0_EFPGA_MATHB_COEF_DATA_14_, MU0_EFPGA_MATHB_COEF_DATA_5_, MU0_EFPGA_MATHB_COEF_DATA_4_, MU0_EFPGA_TPRAM_COEF_W_DATA_31_, MU0_EFPGA_TPRAM_COEF_W_DATA_30_, MU0_EFPGA_MATHB_COEF_DATA_3_, MU0_EFPGA_MATHB_COEF_DATA_2_, MU0_EFPGA_MATHB_COEF_DATA_1_, MU0_EFPGA_MATHB_COEF_DATA_0_, MU0_EFPGA_MATHB_DATAOUT_SEL_1_, MU0_EFPGA_MATHB_DATAOUT_SEL_0_, MU0_EFPGA_TPRAM_COEF_W_MODE_1_, MU0_EFPGA_TPRAM_COEF_W_MODE_0_, MU0_EFPGA_TPRAM_COEF_W_DATA_29_, MU0_EFPGA_TPRAM_COEF_W_DATA_28_, MU0_EFPGA_TPRAM_COEF_W_DATA_19_, MU0_EFPGA_TPRAM_COEF_W_DATA_18_, MU0_EFPGA_TPRAM_COEF_W_DATA_17_, MU0_EFPGA_TPRAM_COEF_W_DATA_16_, MU0_EFPGA_TPRAM_COEF_W_DATA_15_, MU0_EFPGA_TPRAM_COEF_W_DATA_14_, MU0_EFPGA_TPRAM_COEF_W_DATA_13_, MU0_EFPGA_TPRAM_COEF_W_DATA_12_, MU0_EFPGA_TPRAM_COEF_W_DATA_27_, MU0_EFPGA_TPRAM_COEF_W_DATA_26_, MU0_EFPGA_TPRAM_COEF_W_DATA_25_, MU0_EFPGA_TPRAM_COEF_W_DATA_24_, MU0_EFPGA_TPRAM_COEF_W_DATA_23_, MU0_EFPGA_TPRAM_COEF_W_DATA_22_, MU0_EFPGA_TPRAM_COEF_W_DATA_21_, MU0_EFPGA_TPRAM_COEF_W_DATA_20_, MU0_EFPGA_TPRAM_COEF_W_DATA_11_, MU0_EFPGA_TPRAM_COEF_W_DATA_10_, MU0_EFPGA_TPRAM_COEF_W_DATA_1_, MU0_EFPGA_TPRAM_COEF_W_DATA_0_, MU0_EFPGA_TPRAM_COEF_W_DATA_9_, MU0_EFPGA_TPRAM_COEF_W_DATA_8_, MU0_EFPGA_TPRAM_COEF_W_DATA_7_, MU0_EFPGA_TPRAM_COEF_W_DATA_6_, MU0_EFPGA_TPRAM_COEF_W_DATA_5_, MU0_EFPGA_TPRAM_COEF_W_DATA_4_, MU0_EFPGA_TPRAM_COEF_W_DATA_3_, MU0_EFPGA_TPRAM_COEF_W_DATA_2_, MU0_EFPGA_TPRAM_COEF_W_CLK, MU0_EFPGA_TPRAM_COEF_W_ADDR_11_, MU0_EFPGA_TPRAM_COEF_W_ADDR_2_, MU0_EFPGA_TPRAM_COEF_W_ADDR_1_, MU0_EFPGA_TPRAM_COEF_W_ADDR_0_, MU0_EFPGA_TPRAM_COEF_WE, MU0_EFPGA_TPRAM_COEF_WDSEL, MU0_EFPGA_TPRAM_COEF_R_MODE_1_, MU0_EFPGA_TPRAM_COEF_R_MODE_0_, MU0_EFPGA_TPRAM_COEF_R_CLK, MU0_EFPGA_TPRAM_COEF_W_ADDR_10_, MU0_EFPGA_TPRAM_COEF_W_ADDR_9_, MU0_EFPGA_TPRAM_COEF_W_ADDR_8_, MU0_EFPGA_TPRAM_COEF_W_ADDR_7_, MU0_EFPGA_TPRAM_COEF_W_ADDR_6_, MU0_EFPGA_TPRAM_COEF_W_ADDR_5_, MU0_EFPGA_TPRAM_COEF_W_ADDR_4_, MU0_EFPGA_TPRAM_COEF_W_ADDR_3_, MU0_EFPGA_TPRAM_COEF_R_ADDR_11_, MU0_EFPGA_TPRAM_COEF_R_ADDR_10_, MU0_EFPGA_TPRAM_COEF_R_ADDR_1_, MU0_EFPGA_TPRAM_COEF_R_ADDR_0_, MU0_EFPGA_TPRAM_COEF_R_ADDR_9_, MU0_EFPGA_TPRAM_COEF_R_ADDR_8_, MU0_EFPGA_TPRAM_COEF_R_ADDR_7_, MU0_EFPGA_TPRAM_COEF_R_ADDR_6_, MU0_EFPGA_TPRAM_COEF_R_ADDR_5_, MU0_EFPGA_TPRAM_COEF_R_ADDR_4_, MU0_EFPGA_TPRAM_COEF_R_ADDR_3_, MU0_EFPGA_TPRAM_COEF_R_ADDR_2_, MU0_EFPGA_TPRAM_COEF_POWERDN, MU1_EFPGA_TPRAM_OPER_W_MODE_1_, MU1_EFPGA_TPRAM_OPER_W_MODE_0_, MU1_EFPGA_TPRAM_OPER_W_DATA_23_, MU1_EFPGA_TPRAM_OPER_W_DATA_22_, MU1_EFPGA_TPRAM_OPER_W_DATA_31_, MU1_EFPGA_TPRAM_OPER_W_DATA_30_, MU1_EFPGA_TPRAM_OPER_W_DATA_29_, MU1_EFPGA_TPRAM_OPER_W_DATA_28_, MU1_EFPGA_TPRAM_OPER_W_DATA_27_, MU1_EFPGA_TPRAM_OPER_W_DATA_26_, MU1_EFPGA_TPRAM_OPER_W_DATA_25_, MU1_EFPGA_TPRAM_OPER_W_DATA_24_, MU1_EFPGA_TPRAM_OPER_W_DATA_21_, MU1_EFPGA_TPRAM_OPER_W_DATA_20_, MU1_EFPGA_TPRAM_OPER_W_DATA_11_, MU1_EFPGA_TPRAM_OPER_W_DATA_10_, MU1_EFPGA_TPRAM_OPER_W_DATA_9_, MU1_EFPGA_TPRAM_OPER_W_DATA_8_, MU1_EFPGA_TPRAM_OPER_W_DATA_7_, MU1_EFPGA_TPRAM_OPER_W_DATA_6_, MU1_EFPGA_TPRAM_OPER_W_DATA_5_, MU1_EFPGA_TPRAM_OPER_W_DATA_4_, MU1_EFPGA_TPRAM_OPER_W_DATA_19_, MU1_EFPGA_TPRAM_OPER_W_DATA_18_, MU1_EFPGA_TPRAM_OPER_W_DATA_17_, MU1_EFPGA_TPRAM_OPER_W_DATA_16_, MU1_EFPGA_TPRAM_OPER_W_DATA_15_, MU1_EFPGA_TPRAM_OPER_W_DATA_14_, MU1_EFPGA_TPRAM_OPER_W_DATA_13_, MU1_EFPGA_TPRAM_OPER_W_DATA_12_, MU1_EFPGA_TPRAM_OPER_W_DATA_3_, MU1_EFPGA_TPRAM_OPER_W_DATA_2_, MU1_EFPGA_TPRAM_OPER_W_ADDR_6_, MU1_EFPGA_TPRAM_OPER_W_ADDR_5_, MU1_EFPGA_TPRAM_OPER_W_DATA_1_, MU1_EFPGA_TPRAM_OPER_W_DATA_0_, MU1_EFPGA_TPRAM_OPER_W_CLK, MU1_EFPGA_TPRAM_OPER_W_ADDR_11_, MU1_EFPGA_TPRAM_OPER_W_ADDR_10_, MU1_EFPGA_TPRAM_OPER_W_ADDR_9_, MU1_EFPGA_TPRAM_OPER_W_ADDR_8_, MU1_EFPGA_TPRAM_OPER_W_ADDR_7_, MU1_EFPGA_TPRAM_OPER_W_ADDR_4_, MU1_EFPGA_TPRAM_OPER_W_ADDR_3_, MU1_EFPGA_TPRAM_OPER_R_ADDR_11_, MU1_EFPGA_TPRAM_OPER_R_ADDR_10_, MU1_EFPGA_TPRAM_OPER_R_ADDR_9_, MU1_EFPGA_TPRAM_OPER_R_ADDR_8_, MU1_EFPGA_TPRAM_OPER_R_ADDR_7_, MU1_EFPGA_TPRAM_OPER_R_ADDR_6_, MU1_EFPGA_TPRAM_OPER_R_ADDR_5_, MU1_EFPGA_TPRAM_OPER_R_ADDR_4_, MU1_EFPGA_TPRAM_OPER_W_ADDR_2_, MU1_EFPGA_TPRAM_OPER_W_ADDR_1_, MU1_EFPGA_TPRAM_OPER_W_ADDR_0_, MU1_EFPGA_TPRAM_OPER_WE, MU1_EFPGA_TPRAM_OPER_WDSEL, MU1_EFPGA_TPRAM_OPER_R_MODE_1_, MU1_EFPGA_TPRAM_OPER_R_MODE_0_, MU1_EFPGA_TPRAM_OPER_R_CLK, MU1_EFPGA_TPRAM_OPER_R_ADDR_3_, MU1_EFPGA_TPRAM_OPER_R_ADDR_2_, MU1_EFPGA_MATHB_MAC_OUT_SEL_2_, MU1_EFPGA_MATHB_MAC_OUT_SEL_1_, MU1_EFPGA_TPRAM_OPER_R_ADDR_1_, MU1_EFPGA_TPRAM_OPER_R_ADDR_0_, MU1_EFPGA_TPRAM_OPER_POWERDN, MU1_EFPGA2MATHB_CLK, MU1_EFPGA_MATHB_CLK_EN, MU1_EFPGA_MATHB_MAC_OUT_SEL_5_, MU1_EFPGA_MATHB_MAC_OUT_SEL_4_, MU1_EFPGA_MATHB_MAC_OUT_SEL_3_, MU1_EFPGA_MATHB_MAC_OUT_SEL_0_, MU1_EFPGA_MATHB_MAC_ACC_SAT, MU1_EFPGA_MATHB_OPER_DATA_26_, MU1_EFPGA_MATHB_OPER_DATA_25_, MU1_EFPGA_MATHB_OPER_DATA_24_, MU1_EFPGA_MATHB_OPER_DATA_23_, MU1_EFPGA_MATHB_OPER_DATA_22_, MU1_EFPGA_MATHB_OPER_DATA_21_, MU1_EFPGA_MATHB_OPER_DATA_20_, MU1_EFPGA_MATHB_OPER_DATA_19_, MU1_EFPGA_MATHB_MAC_ACC_RND, MU1_EFPGA_MATHB_MAC_ACC_CLEAR, MU1_EFPGA_MATHB_OPER_SEL, MU1_EFPGA_MATHB_OPER_DATA_31_, MU1_EFPGA_MATHB_OPER_DATA_30_, MU1_EFPGA_MATHB_OPER_DATA_29_, MU1_EFPGA_MATHB_OPER_DATA_28_, MU1_EFPGA_MATHB_OPER_DATA_27_, MU1_EFPGA_MATHB_OPER_DATA_18_, MU1_EFPGA_MATHB_OPER_DATA_17_, MU1_EFPGA_MATHB_OPER_DATA_8_, MU1_EFPGA_MATHB_OPER_DATA_7_, MU1_EFPGA_MATHB_OPER_DATA_16_, MU1_EFPGA_MATHB_OPER_DATA_15_, MU1_EFPGA_MATHB_OPER_DATA_14_, MU1_EFPGA_MATHB_OPER_DATA_13_, MU1_EFPGA_MATHB_OPER_DATA_12_, MU1_EFPGA_MATHB_OPER_DATA_11_, MU1_EFPGA_MATHB_OPER_DATA_10_, MU1_EFPGA_MATHB_OPER_DATA_9_, MU1_EFPGA_MATHB_OPER_DATA_6_, MU1_EFPGA_MATHB_OPER_DATA_5_, MU1_EFPGA_MATHB_COEF_DATA_29_, MU1_EFPGA_MATHB_COEF_DATA_28_, MU1_EFPGA_MATHB_COEF_DATA_27_, MU1_EFPGA_MATHB_COEF_DATA_26_, MU1_EFPGA_MATHB_COEF_DATA_25_, MU1_EFPGA_MATHB_COEF_DATA_24_, MU1_EFPGA_MATHB_COEF_DATA_23_, MU1_EFPGA_MATHB_COEF_DATA_22_, MU1_EFPGA_MATHB_OPER_DATA_4_, MU1_EFPGA_MATHB_OPER_DATA_3_, MU1_EFPGA_MATHB_OPER_DATA_2_, MU1_EFPGA_MATHB_OPER_DATA_1_, MU1_EFPGA_MATHB_OPER_DATA_0_, MU1_EFPGA_MATHB_COEF_SEL, MU1_EFPGA_MATHB_COEF_DATA_31_, MU1_EFPGA_MATHB_COEF_DATA_30_, MU1_EFPGA_MATHB_COEF_DATA_21_, MU1_EFPGA_MATHB_COEF_DATA_20_, MU1_EFPGA_MATHB_COEF_DATA_11_, MU1_EFPGA_MATHB_COEF_DATA_10_, MU1_EFPGA_MATHB_COEF_DATA_19_, MU1_EFPGA_MATHB_COEF_DATA_18_, MU1_EFPGA_MATHB_COEF_DATA_17_, MU1_EFPGA_MATHB_COEF_DATA_16_, MU1_EFPGA_MATHB_COEF_DATA_15_, MU1_EFPGA_MATHB_COEF_DATA_14_, MU1_EFPGA_MATHB_COEF_DATA_13_, MU1_EFPGA_MATHB_COEF_DATA_12_, MU1_EFPGA_MATHB_COEF_DATA_9_, MU1_EFPGA_MATHB_COEF_DATA_8_, MU1_EFPGA_MATHB_DATAOUT_SEL_1_, MU1_EFPGA_MATHB_DATAOUT_SEL_0_, MU1_EFPGA_TPRAM_COEF_W_MODE_1_, MU1_EFPGA_TPRAM_COEF_W_MODE_0_, MU1_EFPGA_TPRAM_COEF_W_DATA_31_, MU1_EFPGA_TPRAM_COEF_W_DATA_30_, MU1_EFPGA_TPRAM_COEF_W_DATA_29_, MU1_EFPGA_TPRAM_COEF_W_DATA_28_, MU1_EFPGA_MATHB_COEF_DATA_7_, MU1_EFPGA_MATHB_COEF_DATA_6_, MU1_EFPGA_MATHB_COEF_DATA_5_, MU1_EFPGA_MATHB_COEF_DATA_4_, MU1_EFPGA_MATHB_COEF_DATA_3_, MU1_EFPGA_MATHB_COEF_DATA_2_, MU1_EFPGA_MATHB_COEF_DATA_1_, MU1_EFPGA_MATHB_COEF_DATA_0_, MU1_EFPGA_TPRAM_COEF_W_DATA_27_, MU1_EFPGA_TPRAM_COEF_W_DATA_26_, MU1_EFPGA_TPRAM_COEF_W_DATA_17_, MU1_EFPGA_TPRAM_COEF_W_DATA_16_, MU1_EFPGA_TPRAM_COEF_W_DATA_25_, MU1_EFPGA_TPRAM_COEF_W_DATA_24_, MU1_EFPGA_TPRAM_COEF_W_DATA_23_, MU1_EFPGA_TPRAM_COEF_W_DATA_22_, MU1_EFPGA_TPRAM_COEF_W_DATA_21_, MU1_EFPGA_TPRAM_COEF_W_DATA_20_, MU1_EFPGA_TPRAM_COEF_W_DATA_19_, MU1_EFPGA_TPRAM_COEF_W_DATA_18_, MU1_EFPGA_TPRAM_COEF_W_DATA_15_, MU1_EFPGA_TPRAM_COEF_W_DATA_14_, MU1_EFPGA_TPRAM_COEF_W_DATA_5_, MU1_EFPGA_TPRAM_COEF_W_DATA_4_, MU1_EFPGA_TPRAM_COEF_W_DATA_3_, MU1_EFPGA_TPRAM_COEF_W_DATA_2_, MU1_EFPGA_TPRAM_COEF_W_DATA_1_, MU1_EFPGA_TPRAM_COEF_W_DATA_0_, MU1_EFPGA_TPRAM_COEF_W_CLK, MU1_EFPGA_TPRAM_COEF_W_ADDR_11_, MU1_EFPGA_TPRAM_COEF_W_DATA_13_, MU1_EFPGA_TPRAM_COEF_W_DATA_12_, MU1_EFPGA_TPRAM_COEF_W_DATA_11_, MU1_EFPGA_TPRAM_COEF_W_DATA_10_, MU1_EFPGA_TPRAM_COEF_W_DATA_9_, MU1_EFPGA_TPRAM_COEF_W_DATA_8_, MU1_EFPGA_TPRAM_COEF_W_DATA_7_, MU1_EFPGA_TPRAM_COEF_W_DATA_6_, MU1_EFPGA_TPRAM_COEF_W_ADDR_10_, MU1_EFPGA_TPRAM_COEF_W_ADDR_9_, MU1_EFPGA_TPRAM_COEF_W_ADDR_0_, MU1_EFPGA_TPRAM_COEF_WE, MU1_EFPGA_TPRAM_COEF_W_ADDR_8_, MU1_EFPGA_TPRAM_COEF_W_ADDR_7_, MU1_EFPGA_TPRAM_COEF_W_ADDR_6_, MU1_EFPGA_TPRAM_COEF_W_ADDR_5_, MU1_EFPGA_TPRAM_COEF_W_ADDR_4_, MU1_EFPGA_TPRAM_COEF_W_ADDR_3_, MU1_EFPGA_TPRAM_COEF_W_ADDR_2_, MU1_EFPGA_TPRAM_COEF_W_ADDR_1_, MU0_EFPGA_TPRAM_OPER_W_DATA_25_, MU0_EFPGA_TPRAM_OPER_W_DATA_24_, MU0_EFPGA_TPRAM_OPER_W_DATA_23_, MU0_EFPGA_TPRAM_OPER_W_DATA_22_, MU0_EFPGA_TPRAM_OPER_W_DATA_21_, MU0_EFPGA_TPRAM_OPER_W_DATA_20_, MU0_EFPGA_TPRAM_OPER_W_DATA_19_, MU0_EFPGA_TPRAM_OPER_W_DATA_18_, MU0_EFPGA_TPRAM_OPER_W_MODE_1_, MU0_EFPGA_TPRAM_OPER_W_MODE_0_, MU0_EFPGA_TPRAM_OPER_W_DATA_31_, MU0_EFPGA_TPRAM_OPER_W_DATA_30_, MU0_EFPGA_TPRAM_OPER_W_DATA_29_, MU0_EFPGA_TPRAM_OPER_W_DATA_28_, MU0_EFPGA_TPRAM_OPER_W_DATA_27_, MU0_EFPGA_TPRAM_OPER_W_DATA_26_, MU1_EFPGA_TPRAM_COEF_WDSEL, MU1_EFPGA_TPRAM_COEF_R_MODE_1_, MU1_EFPGA_TPRAM_COEF_R_ADDR_5_, MU1_EFPGA_TPRAM_COEF_R_ADDR_4_, MU1_EFPGA_TPRAM_COEF_R_ADDR_3_, MU1_EFPGA_TPRAM_COEF_R_ADDR_2_, MU1_EFPGA_TPRAM_COEF_R_ADDR_1_, MU1_EFPGA_TPRAM_COEF_R_ADDR_0_, MU1_EFPGA_TPRAM_COEF_POWERDN, MU1_EFPGA_TPRAM_COEF_R_MODE_0_, MU1_EFPGA_TPRAM_COEF_R_CLK, MU1_EFPGA_TPRAM_COEF_R_ADDR_11_, MU1_EFPGA_TPRAM_COEF_R_ADDR_10_, MU1_EFPGA_TPRAM_COEF_R_ADDR_9_, MU1_EFPGA_TPRAM_COEF_R_ADDR_8_, MU1_EFPGA_TPRAM_COEF_R_ADDR_7_, MU1_EFPGA_TPRAM_COEF_R_ADDR_6_, MU0_EFPGA_TPRAM_OPER_W_DATA_17_, MU0_EFPGA_TPRAM_OPER_W_DATA_16_, MU0_EFPGA_TPRAM_OPER_W_DATA_7_, MU0_EFPGA_TPRAM_OPER_W_DATA_6_, MU0_EFPGA_TPRAM_OPER_W_DATA_15_, MU0_EFPGA_TPRAM_OPER_W_DATA_14_, MU0_EFPGA_TPRAM_OPER_W_DATA_13_, MU0_EFPGA_TPRAM_OPER_W_DATA_12_, MU0_EFPGA_TPRAM_OPER_W_DATA_11_, MU0_EFPGA_TPRAM_OPER_W_DATA_10_, MU0_EFPGA_TPRAM_OPER_W_DATA_9_, MU0_EFPGA_TPRAM_OPER_W_DATA_8_, MU0_EFPGA_TPRAM_OPER_W_DATA_5_, MU0_EFPGA_TPRAM_OPER_W_DATA_4_, MU0_EFPGA_TPRAM_OPER_W_ADDR_8_, MU0_EFPGA_TPRAM_OPER_W_ADDR_7_, MU0_EFPGA_TPRAM_OPER_W_ADDR_6_, MU0_EFPGA_TPRAM_OPER_W_ADDR_5_, MU0_EFPGA_TPRAM_OPER_W_ADDR_4_, MU0_EFPGA_TPRAM_OPER_W_ADDR_3_, MU0_EFPGA_TPRAM_OPER_W_ADDR_2_, MU0_EFPGA_TPRAM_OPER_W_ADDR_1_, MU0_EFPGA_TPRAM_OPER_W_DATA_3_, MU0_EFPGA_TPRAM_OPER_W_DATA_2_, MU0_EFPGA_TPRAM_OPER_W_DATA_1_, MU0_EFPGA_TPRAM_OPER_W_DATA_0_, MU0_EFPGA_TPRAM_OPER_W_CLK, MU0_EFPGA_TPRAM_OPER_W_ADDR_11_, MU0_EFPGA_TPRAM_OPER_W_ADDR_10_, MU0_EFPGA_TPRAM_OPER_W_ADDR_9_, MU0_EFPGA_TPRAM_OPER_W_ADDR_0_, MU0_EFPGA_TPRAM_OPER_WE, MU0_EFPGA_TPRAM_OPER_R_ADDR_7_, MU0_EFPGA_TPRAM_OPER_R_ADDR_6_, MU0_EFPGA_TPRAM_OPER_WDSEL, MU0_EFPGA_TPRAM_OPER_R_MODE_1_, MU0_EFPGA_TPRAM_OPER_R_MODE_0_, MU0_EFPGA_TPRAM_OPER_R_CLK, MU0_EFPGA_TPRAM_OPER_R_ADDR_11_, MU0_EFPGA_TPRAM_OPER_R_ADDR_10_, MU0_EFPGA_TPRAM_OPER_R_ADDR_9_, MU0_EFPGA_TPRAM_OPER_R_ADDR_8_, MU0_EFPGA_TPRAM_OPER_R_ADDR_5_, MU0_EFPGA_TPRAM_OPER_R_ADDR_4_, MU0_EFPGA_MATHB_MAC_OUT_SEL_4_, MU0_EFPGA_MATHB_MAC_OUT_SEL_3_, MU0_EFPGA_MATHB_MAC_OUT_SEL_2_, MU0_EFPGA_MATHB_MAC_OUT_SEL_1_, MU0_EFPGA_MATHB_MAC_OUT_SEL_0_, MU0_EFPGA_MATHB_MAC_ACC_SAT, MU0_EFPGA_MATHB_MAC_ACC_RND, MU0_EFPGA_MATHB_MAC_ACC_CLEAR, MU0_EFPGA_TPRAM_OPER_R_ADDR_3_, MU0_EFPGA_TPRAM_OPER_R_ADDR_2_, MU0_EFPGA_TPRAM_OPER_R_ADDR_1_, MU0_EFPGA_TPRAM_OPER_R_ADDR_0_, MU0_EFPGA_TPRAM_OPER_POWERDN, MU0_EFPGA2MATHB_CLK, MU0_EFPGA_MATHB_CLK_EN, MU0_EFPGA_MATHB_MAC_OUT_SEL_5_, MU0_EFPGA_MATHB_OPER_SEL, MU0_EFPGA_MATHB_OPER_DATA_31_, MU0_EFPGA_MATHB_OPER_DATA_22_, MU0_EFPGA_MATHB_OPER_DATA_21_, MU0_EFPGA_MATHB_OPER_DATA_30_, MU0_EFPGA_MATHB_OPER_DATA_29_, MU0_EFPGA_MATHB_OPER_DATA_28_, MU0_EFPGA_MATHB_OPER_DATA_27_, MU0_EFPGA_MATHB_OPER_DATA_26_, MU0_EFPGA_MATHB_OPER_DATA_25_, MU0_EFPGA_MATHB_OPER_DATA_24_, MU0_EFPGA_MATHB_OPER_DATA_23_, MU0_EFPGA_MATHB_OPER_DATA_20_, MU0_EFPGA_MATHB_OPER_DATA_19_, MU0_EFPGA_MATHB_OPER_DATA_10_, MU0_EFPGA_MATHB_OPER_DATA_9_, MU0_EFPGA_MATHB_OPER_DATA_8_, MU0_EFPGA_MATHB_OPER_DATA_7_, MU0_EFPGA_MATHB_OPER_DATA_6_, MU0_EFPGA_MATHB_OPER_DATA_5_, MU0_EFPGA_MATHB_OPER_DATA_4_, MU0_EFPGA_MATHB_OPER_DATA_3_, MU0_EFPGA_MATHB_OPER_DATA_18_, MU0_EFPGA_MATHB_OPER_DATA_17_, MU0_EFPGA_MATHB_OPER_DATA_16_, MU0_EFPGA_MATHB_OPER_DATA_15_, MU0_EFPGA_MATHB_OPER_DATA_14_, MU0_EFPGA_MATHB_OPER_DATA_13_, MU0_EFPGA_MATHB_OPER_DATA_12_, MU0_EFPGA_MATHB_OPER_DATA_11_, MU0_EFPGA_MATHB_OPER_DATA_2_, MU0_EFPGA_MATHB_OPER_DATA_1_, MU0_EFPGA_MATHB_COEF_DATA_25_, MU0_EFPGA_MATHB_COEF_DATA_24_, MU0_EFPGA_MATHB_OPER_DATA_0_, MU0_EFPGA_MATHB_COEF_SEL, MU0_EFPGA_MATHB_COEF_DATA_31_, MU0_EFPGA_MATHB_COEF_DATA_30_, MU0_EFPGA_MATHB_COEF_DATA_29_, MU0_EFPGA_MATHB_COEF_DATA_28_, MU0_EFPGA_MATHB_COEF_DATA_27_, MU0_EFPGA_MATHB_COEF_DATA_26_, MU1_EFPGA_MATHB_TC_defPin, MU1_EFPGA_MATHB_OPER_defPin_1_, MU1_EFPGA_MATHB_OPER_defPin_0_, MU1_EFPGA_MATHB_COEF_defPin_1_, MU1_EFPGA_MATHB_COEF_defPin_0_, MU0_EFPGA_MATHB_TC_defPin, MU0_EFPGA_MATHB_OPER_defPin_1_, MU0_EFPGA_MATHB_OPER_defPin_0_, MU0_EFPGA_MATHB_COEF_defPin_1_, MU0_EFPGA_MATHB_COEF_defPin_0_, BL_DOUT_0_, BL_DOUT_10_, BL_DOUT_11_, BL_DOUT_12_, BL_DOUT_13_, BL_DOUT_14_, BL_DOUT_15_, BL_DOUT_16_, BL_DOUT_17_, BL_DOUT_18_, BL_DOUT_19_, BL_DOUT_1_, BL_DOUT_20_, BL_DOUT_21_, BL_DOUT_22_, BL_DOUT_23_, BL_DOUT_24_, BL_DOUT_25_, BL_DOUT_26_, BL_DOUT_27_, BL_DOUT_28_, BL_DOUT_29_, BL_DOUT_2_, BL_DOUT_30_, BL_DOUT_31_, BL_DOUT_3_, BL_DOUT_4_, BL_DOUT_5_, BL_DOUT_6_, BL_DOUT_7_, BL_DOUT_8_, BL_DOUT_9_, FB_SPE_OUT_0_, FB_SPE_OUT_1_, FB_SPE_OUT_2_, FB_SPE_OUT_3_, PARALLEL_CFG;

QL_eFPGA_ArcticPro2_32X32_GF_22_QL_eFPGA myDeviceInstance_QL_eFPGA_ArcticPro2_32X32_GF_22_QL_eFPGA (
.A2F_CLK0(CLK0),
.A2F_CLK1(CLK1),
.A2F_CLK2(CLK2),
.A2F_CLK3(CLK3),
.A2F_CLK4(CLK4),
.A2F_CLK5(CLK5),
.A2F_B_10_0(supplyBus[0]),
.A2F_B_10_1(supplyBus[1]),
.A2F_B_10_2(supplyBus[2]),
.A2F_B_10_3(supplyBus[3]),
.A2F_B_10_4(supplyBus[4]),
.A2F_B_10_5(supplyBus[5]),
.A2F_B_10_6(supplyBus[6]),
.A2F_B_10_7(supplyBus[7]),
.A2F_B_11_0(supplyBus[8]),
.A2F_B_11_1(supplyBus[9]),
.A2F_B_11_2(supplyBus[10]),
.A2F_B_11_3(supplyBus[11]),
.A2F_B_11_4(supplyBus[12]),
.A2F_B_11_5(supplyBus[13]),
.A2F_B_12_0(supplyBus[14]),
.A2F_B_12_1(supplyBus[15]),
.A2F_B_12_2(supplyBus[16]),
.A2F_B_12_3(supplyBus[17]),
.A2F_B_12_4(supplyBus[18]),
.A2F_B_12_5(supplyBus[19]),
.A2F_B_12_6(supplyBus[20]),
.A2F_B_12_7(supplyBus[21]),
.A2F_B_13_0(supplyBus[22]),
.A2F_B_13_1(supplyBus[23]),
.A2F_B_13_2(supplyBus[24]),
.A2F_B_13_3(supplyBus[25]),
.A2F_B_13_4(supplyBus[26]),
.A2F_B_13_5(supplyBus[27]),
.A2F_B_14_0(supplyBus[28]),
.A2F_B_14_1(supplyBus[29]),
.A2F_B_14_2(supplyBus[30]),
.A2F_B_14_3(supplyBus[31]),
.A2F_B_14_4(supplyBus[32]),
.A2F_B_14_5(supplyBus[33]),
.A2F_B_14_6(supplyBus[34]),
.A2F_B_14_7(supplyBus[35]),
.A2F_B_15_0(supplyBus[36]),
.A2F_B_15_1(supplyBus[37]),
.A2F_B_15_2(supplyBus[38]),
.A2F_B_15_3(supplyBus[39]),
.A2F_B_15_4(supplyBus[40]),
.A2F_B_15_5(supplyBus[41]),
.A2F_B_16_0(fpgaio_data_0_i),
.A2F_B_16_1(fpgaio_data_1_i),
.A2F_B_16_2(fpgaio_data_2_i),
.A2F_B_16_3(fpgaio_data_3_i),
.A2F_B_16_4(supplyBus[42]),
.A2F_B_16_5(supplyBus[43]),
.A2F_B_16_6(supplyBus[44]),
.A2F_B_16_7(supplyBus[45]),
.A2F_B_17_0(fpgaio_data_4_i),
.A2F_B_17_1(fpgaio_data_5_i),
.A2F_B_17_2(fpgaio_data_6_i),
.A2F_B_17_3(fpgaio_data_7_i),
.A2F_B_17_4(supplyBus[46]),
.A2F_B_17_5(supplyBus[47]),
.A2F_B_18_0(supplyBus[48]),
.A2F_B_18_1(supplyBus[49]),
.A2F_B_18_2(supplyBus[50]),
.A2F_B_18_3(supplyBus[51]),
.A2F_B_18_4(supplyBus[52]),
.A2F_B_18_5(supplyBus[53]),
.A2F_B_18_6(supplyBus[54]),
.A2F_B_18_7(supplyBus[55]),
.A2F_B_19_0(supplyBus[56]),
.A2F_B_19_1(supplyBus[57]),
.A2F_B_19_2(supplyBus[58]),
.A2F_B_19_3(supplyBus[59]),
.A2F_B_19_4(supplyBus[60]),
.A2F_B_19_5(supplyBus[61]),
.A2F_B_1_0(supplyBus[62]),
.A2F_B_1_1(supplyBus[63]),
.A2F_B_1_2(supplyBus[64]),
.A2F_B_1_3(supplyBus[65]),
.A2F_B_1_4(supplyBus[66]),
.A2F_B_1_5(supplyBus[67]),
.A2F_B_20_0(supplyBus[68]),
.A2F_B_20_1(supplyBus[69]),
.A2F_B_20_2(supplyBus[70]),
.A2F_B_20_3(supplyBus[71]),
.A2F_B_20_4(supplyBus[72]),
.A2F_B_20_5(supplyBus[73]),
.A2F_B_20_6(supplyBus[74]),
.A2F_B_20_7(supplyBus[75]),
.A2F_B_21_0(supplyBus[76]),
.A2F_B_21_1(supplyBus[77]),
.A2F_B_21_2(supplyBus[78]),
.A2F_B_21_3(supplyBus[79]),
.A2F_B_21_4(supplyBus[80]),
.A2F_B_21_5(supplyBus[81]),
.A2F_B_22_0(supplyBus[82]),
.A2F_B_22_1(supplyBus[83]),
.A2F_B_22_2(supplyBus[84]),
.A2F_B_22_3(supplyBus[85]),
.A2F_B_22_4(supplyBus[86]),
.A2F_B_22_5(supplyBus[87]),
.A2F_B_22_6(supplyBus[88]),
.A2F_B_22_7(supplyBus[89]),
.A2F_B_23_0(supplyBus[90]),
.A2F_B_23_1(supplyBus[91]),
.A2F_B_23_2(supplyBus[92]),
.A2F_B_23_3(supplyBus[93]),
.A2F_B_23_4(supplyBus[94]),
.A2F_B_23_5(supplyBus[95]),
.A2F_B_24_0(supplyBus[96]),
.A2F_B_24_1(supplyBus[97]),
.A2F_B_24_2(supplyBus[98]),
.A2F_B_24_3(supplyBus[99]),
.A2F_B_24_4(supplyBus[100]),
.A2F_B_24_5(supplyBus[101]),
.A2F_B_24_6(supplyBus[102]),
.A2F_B_24_7(supplyBus[103]),
.A2F_B_25_0(supplyBus[104]),
.A2F_B_25_1(supplyBus[105]),
.A2F_B_25_2(supplyBus[106]),
.A2F_B_25_3(supplyBus[107]),
.A2F_B_25_4(supplyBus[108]),
.A2F_B_25_5(supplyBus[109]),
.A2F_B_26_0(supplyBus[110]),
.A2F_B_26_1(supplyBus[111]),
.A2F_B_26_2(supplyBus[112]),
.A2F_B_26_3(supplyBus[113]),
.A2F_B_26_4(supplyBus[114]),
.A2F_B_26_5(supplyBus[115]),
.A2F_B_26_6(supplyBus[116]),
.A2F_B_26_7(supplyBus[117]),
.A2F_B_27_0(supplyBus[118]),
.A2F_B_27_1(supplyBus[119]),
.A2F_B_27_2(supplyBus[120]),
.A2F_B_27_3(supplyBus[121]),
.A2F_B_27_4(supplyBus[122]),
.A2F_B_27_5(supplyBus[123]),
.A2F_B_28_0(supplyBus[124]),
.A2F_B_28_1(supplyBus[125]),
.A2F_B_28_2(supplyBus[126]),
.A2F_B_28_3(supplyBus[127]),
.A2F_B_28_4(supplyBus[128]),
.A2F_B_28_5(supplyBus[129]),
.A2F_B_28_6(supplyBus[130]),
.A2F_B_28_7(supplyBus[131]),
.A2F_B_29_0(supplyBus[132]),
.A2F_B_29_1(supplyBus[133]),
.A2F_B_29_2(supplyBus[134]),
.A2F_B_29_3(supplyBus[135]),
.A2F_B_29_4(supplyBus[136]),
.A2F_B_29_5(supplyBus[137]),
.A2F_B_2_0(supplyBus[138]),
.A2F_B_2_1(supplyBus[139]),
.A2F_B_2_2(supplyBus[140]),
.A2F_B_2_3(supplyBus[141]),
.A2F_B_2_4(supplyBus[142]),
.A2F_B_2_5(supplyBus[143]),
.A2F_B_2_6(supplyBus[144]),
.A2F_B_2_7(supplyBus[145]),
.A2F_B_30_0(supplyBus[146]),
.A2F_B_30_1(supplyBus[147]),
.A2F_B_30_2(supplyBus[148]),
.A2F_B_30_3(supplyBus[149]),
.A2F_B_30_4(supplyBus[150]),
.A2F_B_30_5(supplyBus[151]),
.A2F_B_30_6(supplyBus[152]),
.A2F_B_30_7(supplyBus[153]),
.A2F_B_31_0(supplyBus[154]),
.A2F_B_31_1(supplyBus[155]),
.A2F_B_31_2(supplyBus[156]),
.A2F_B_31_3(supplyBus[157]),
.A2F_B_31_4(supplyBus[158]),
.A2F_B_31_5(supplyBus[159]),
.A2F_B_32_0(supplyBus[160]),
.A2F_B_32_1(supplyBus[161]),
.A2F_B_32_2(supplyBus[162]),
.A2F_B_32_3(supplyBus[163]),
.A2F_B_32_4(supplyBus[164]),
.A2F_B_32_5(supplyBus[165]),
.A2F_B_32_6(supplyBus[166]),
.A2F_B_32_7(supplyBus[167]),
.A2F_B_3_0(supplyBus[168]),
.A2F_B_3_1(supplyBus[169]),
.A2F_B_3_2(supplyBus[170]),
.A2F_B_3_3(supplyBus[171]),
.A2F_B_3_4(supplyBus[172]),
.A2F_B_3_5(supplyBus[173]),
.A2F_B_4_0(supplyBus[174]),
.A2F_B_4_1(supplyBus[175]),
.A2F_B_4_2(supplyBus[176]),
.A2F_B_4_3(supplyBus[177]),
.A2F_B_4_4(supplyBus[178]),
.A2F_B_4_5(supplyBus[179]),
.A2F_B_4_6(supplyBus[180]),
.A2F_B_4_7(supplyBus[181]),
.A2F_B_5_0(supplyBus[182]),
.A2F_B_5_1(supplyBus[183]),
.A2F_B_5_2(supplyBus[184]),
.A2F_B_5_3(supplyBus[185]),
.A2F_B_5_4(supplyBus[186]),
.A2F_B_5_5(supplyBus[187]),
.A2F_B_6_0(supplyBus[188]),
.A2F_B_6_1(supplyBus[189]),
.A2F_B_6_2(supplyBus[190]),
.A2F_B_6_3(supplyBus[191]),
.A2F_B_6_4(supplyBus[192]),
.A2F_B_6_5(supplyBus[193]),
.A2F_B_6_6(supplyBus[194]),
.A2F_B_6_7(supplyBus[195]),
.A2F_B_7_0(supplyBus[196]),
.A2F_B_7_1(supplyBus[197]),
.A2F_B_7_2(supplyBus[198]),
.A2F_B_7_3(supplyBus[199]),
.A2F_B_7_4(supplyBus[200]),
.A2F_B_7_5(supplyBus[201]),
.A2F_B_8_0(supplyBus[202]),
.A2F_B_8_1(supplyBus[203]),
.A2F_B_8_2(supplyBus[204]),
.A2F_B_8_3(supplyBus[205]),
.A2F_B_8_4(supplyBus[206]),
.A2F_B_8_5(supplyBus[207]),
.A2F_B_8_6(supplyBus[208]),
.A2F_B_8_7(supplyBus[209]),
.A2F_B_9_0(supplyBus[210]),
.A2F_B_9_1(supplyBus[211]),
.A2F_B_9_2(supplyBus[212]),
.A2F_B_9_3(supplyBus[213]),
.A2F_B_9_4(supplyBus[214]),
.A2F_B_9_5(supplyBus[215]),
.A2F_L_10_0(udma_cfg_data_8_i),
.A2F_L_10_1(udma_cfg_data_9_i),
.A2F_L_10_2(udma_cfg_data_10_i),
.A2F_L_10_3(udma_cfg_data_11_i),
.A2F_L_10_4(udma_cfg_data_12_i),
.A2F_L_10_5(udma_cfg_data_13_i),
.A2F_L_10_6(udma_cfg_data_14_i),
.A2F_L_10_7(udma_cfg_data_15_i),
.A2F_L_11_0(udma_cfg_data_2_i),
.A2F_L_11_1(udma_cfg_data_3_i),
.A2F_L_11_2(udma_cfg_data_4_i),
.A2F_L_11_3(udma_cfg_data_5_i),
.A2F_L_11_4(udma_cfg_data_6_i),
.A2F_L_11_5(udma_cfg_data_7_i),
.A2F_L_12_0(udma_tx_lin_data_27_i),
.A2F_L_12_1(udma_tx_lin_data_28_i),
.A2F_L_12_2(udma_tx_lin_data_29_i),
.A2F_L_12_3(udma_tx_lin_data_30_i),
.A2F_L_12_4(udma_tx_lin_data_31_i),
.A2F_L_12_5(udma_rx_lin_ready_i),
.A2F_L_12_6(udma_cfg_data_0_i),
.A2F_L_12_7(udma_cfg_data_1_i),
.A2F_L_13_0(udma_tx_lin_data_21_i),
.A2F_L_13_1(udma_tx_lin_data_22_i),
.A2F_L_13_2(udma_tx_lin_data_23_i),
.A2F_L_13_3(udma_tx_lin_data_24_i),
.A2F_L_13_4(udma_tx_lin_data_25_i),
.A2F_L_13_5(udma_tx_lin_data_26_i),
.A2F_L_14_0(udma_tx_lin_data_13_i),
.A2F_L_14_1(udma_tx_lin_data_14_i),
.A2F_L_14_2(udma_tx_lin_data_15_i),
.A2F_L_14_3(udma_tx_lin_data_16_i),
.A2F_L_14_4(udma_tx_lin_data_17_i),
.A2F_L_14_5(udma_tx_lin_data_18_i),
.A2F_L_14_6(udma_tx_lin_data_19_i),
.A2F_L_14_7(udma_tx_lin_data_20_i),
.A2F_L_15_0(udma_tx_lin_data_7_i),
.A2F_L_15_1(udma_tx_lin_data_8_i),
.A2F_L_15_2(udma_tx_lin_data_9_i),
.A2F_L_15_3(udma_tx_lin_data_10_i),
.A2F_L_15_4(udma_tx_lin_data_11_i),
.A2F_L_15_5(udma_tx_lin_data_12_i),
.A2F_L_16_0(udma_tx_lin_valid_i),
.A2F_L_16_1(udma_tx_lin_data_0_i),
.A2F_L_16_2(udma_tx_lin_data_1_i),
.A2F_L_16_3(udma_tx_lin_data_2_i),
.A2F_L_16_4(udma_tx_lin_data_3_i),
.A2F_L_16_5(udma_tx_lin_data_4_i),
.A2F_L_16_6(udma_tx_lin_data_5_i),
.A2F_L_16_7(udma_tx_lin_data_6_i),
.A2F_L_17_0(apb_hwce_pwdata_0_i),
.A2F_L_17_1(apb_hwce_pwdata_1_i),
.A2F_L_17_2(apb_hwce_pwdata_2_i),
.A2F_L_17_3(apb_hwce_pwdata_3_i),
.A2F_L_17_4(apb_hwce_pwdata_4_i),
.A2F_L_17_5(apb_hwce_pwdata_5_i),
.A2F_L_18_0(apb_hwce_pwdata_6_i),
.A2F_L_18_1(apb_hwce_pwdata_7_i),
.A2F_L_18_2(apb_hwce_pwdata_8_i),
.A2F_L_18_3(apb_hwce_pwdata_9_i),
.A2F_L_18_4(apb_hwce_pwdata_10_i),
.A2F_L_18_5(apb_hwce_pwdata_11_i),
.A2F_L_18_6(apb_hwce_pwdata_12_i),
.A2F_L_18_7(apb_hwce_pwdata_13_i),
.A2F_L_19_0(apb_hwce_pwdata_14_i),
.A2F_L_19_1(apb_hwce_pwdata_15_i),
.A2F_L_19_2(apb_hwce_pwdata_16_i),
.A2F_L_19_3(apb_hwce_pwdata_17_i),
.A2F_L_19_4(apb_hwce_pwdata_18_i),
.A2F_L_19_5(apb_hwce_pwdata_19_i),
.A2F_L_1_0(supplyBus[216]),
.A2F_L_1_1(supplyBus[217]),
.A2F_L_1_2(supplyBus[218]),
.A2F_L_1_3(supplyBus[219]),
.A2F_L_1_4(supplyBus[220]),
.A2F_L_1_5(supplyBus[221]),
.A2F_L_20_0(apb_hwce_pwdata_20_i),
.A2F_L_20_1(apb_hwce_pwdata_21_i),
.A2F_L_20_2(apb_hwce_pwdata_22_i),
.A2F_L_20_3(apb_hwce_pwdata_23_i),
.A2F_L_20_4(apb_hwce_pwdata_24_i),
.A2F_L_20_5(apb_hwce_pwdata_25_i),
.A2F_L_20_6(apb_hwce_pwdata_26_i),
.A2F_L_20_7(apb_hwce_pwdata_27_i),
.A2F_L_21_0(apb_hwce_pwdata_28_i),
.A2F_L_21_1(apb_hwce_pwdata_29_i),
.A2F_L_21_2(apb_hwce_pwdata_30_i),
.A2F_L_21_3(apb_hwce_pwdata_31_i),
.A2F_L_21_4(apb_hwce_addr_0_i),
.A2F_L_21_5(apb_hwce_addr_1_i),
.A2F_L_22_0(apb_hwce_addr_2_i),
.A2F_L_22_1(apb_hwce_addr_3_i),
.A2F_L_22_2(apb_hwce_addr_4_i),
.A2F_L_22_3(apb_hwce_addr_5_i),
.A2F_L_22_4(apb_hwce_addr_6_i),
.A2F_L_22_5(apb_hwce_enable_i),
.A2F_L_22_6(apb_hwce_psel_i),
.A2F_L_22_7(apb_hwce_pstrb_i),
.A2F_L_23_0(apb_hwce_pwrite_i),
.A2F_L_23_1(fpgaio_data_28_i),
.A2F_L_23_2(fpgaio_data_29_i),
.A2F_L_23_3(fpgaio_data_30_i),
.A2F_L_23_4(fpgaio_data_31_i),
.A2F_L_23_5(fpgaio_data_32_i),
.A2F_L_24_0(fpgaio_data_33_i),
.A2F_L_24_1(fpgaio_data_34_i),
.A2F_L_24_2(fpgaio_data_35_i),
.A2F_L_24_3(fpgaio_data_36_i),
.A2F_L_24_4(fpgaio_data_37_i),
.A2F_L_24_5(fpgaio_data_38_i),
.A2F_L_24_6(fpgaio_data_39_i),
.A2F_L_24_7(fpgaio_data_40_i),
.A2F_L_25_0(fpgaio_data_41_i),
.A2F_L_25_1(fpgaio_data_42_i),
.A2F_L_25_2(RESET_LB),
.A2F_L_25_3(supplyBus[222]),
.A2F_L_25_4(supplyBus[223]),
.A2F_L_25_5(supplyBus[224]),
.A2F_L_26_0(supplyBus[225]),
.A2F_L_26_1(supplyBus[226]),
.A2F_L_26_2(supplyBus[227]),
.A2F_L_26_3(supplyBus[228]),
.A2F_L_26_4(supplyBus[229]),
.A2F_L_26_5(supplyBus[230]),
.A2F_L_26_6(supplyBus[231]),
.A2F_L_26_7(supplyBus[232]),
.A2F_L_27_0(supplyBus[233]),
.A2F_L_27_1(supplyBus[234]),
.A2F_L_27_2(supplyBus[235]),
.A2F_L_27_3(supplyBus[236]),
.A2F_L_27_4(supplyBus[237]),
.A2F_L_27_5(supplyBus[238]),
.A2F_L_28_0(supplyBus[239]),
.A2F_L_28_1(supplyBus[240]),
.A2F_L_28_2(supplyBus[241]),
.A2F_L_28_3(supplyBus[242]),
.A2F_L_28_4(supplyBus[243]),
.A2F_L_28_5(supplyBus[244]),
.A2F_L_28_6(supplyBus[245]),
.A2F_L_28_7(supplyBus[246]),
.A2F_L_29_0(supplyBus[247]),
.A2F_L_29_1(supplyBus[248]),
.A2F_L_29_2(supplyBus[249]),
.A2F_L_29_3(supplyBus[250]),
.A2F_L_29_4(supplyBus[251]),
.A2F_L_29_5(supplyBus[252]),
.A2F_L_2_0(supplyBus[253]),
.A2F_L_2_1(supplyBus[254]),
.A2F_L_2_2(supplyBus[255]),
.A2F_L_2_3(supplyBus[256]),
.A2F_L_2_4(supplyBus[257]),
.A2F_L_2_5(supplyBus[258]),
.A2F_L_2_6(supplyBus[259]),
.A2F_L_2_7(supplyBus[260]),
.A2F_L_30_0(supplyBus[261]),
.A2F_L_30_1(supplyBus[262]),
.A2F_L_30_2(supplyBus[263]),
.A2F_L_30_3(supplyBus[264]),
.A2F_L_30_4(supplyBus[265]),
.A2F_L_30_5(supplyBus[266]),
.A2F_L_30_6(supplyBus[267]),
.A2F_L_30_7(supplyBus[268]),
.A2F_L_31_0(supplyBus[269]),
.A2F_L_31_1(supplyBus[270]),
.A2F_L_31_2(supplyBus[271]),
.A2F_L_31_3(supplyBus[272]),
.A2F_L_31_4(supplyBus[273]),
.A2F_L_31_5(supplyBus[274]),
.A2F_L_32_0(supplyBus[275]),
.A2F_L_32_1(supplyBus[276]),
.A2F_L_32_2(supplyBus[277]),
.A2F_L_32_3(supplyBus[278]),
.A2F_L_32_4(supplyBus[279]),
.A2F_L_32_5(supplyBus[280]),
.A2F_L_32_6(supplyBus[281]),
.A2F_L_32_7(supplyBus[282]),
.A2F_L_3_0(supplyBus[283]),
.A2F_L_3_1(supplyBus[284]),
.A2F_L_3_2(supplyBus[285]),
.A2F_L_3_3(supplyBus[286]),
.A2F_L_3_4(supplyBus[287]),
.A2F_L_3_5(supplyBus[288]),
.A2F_L_4_0(supplyBus[289]),
.A2F_L_4_1(supplyBus[290]),
.A2F_L_4_2(supplyBus[291]),
.A2F_L_4_3(supplyBus[292]),
.A2F_L_4_4(supplyBus[293]),
.A2F_L_4_5(supplyBus[294]),
.A2F_L_4_6(supplyBus[295]),
.A2F_L_4_7(supplyBus[296]),
.A2F_L_5_0(RESET_LT),
.A2F_L_5_1(supplyBus[297]),
.A2F_L_5_2(supplyBus[298]),
.A2F_L_5_3(supplyBus[299]),
.A2F_L_5_4(supplyBus[300]),
.A2F_L_5_5(supplyBus[301]),
.A2F_L_6_0(fpgaio_data_20_i),
.A2F_L_6_1(fpgaio_data_21_i),
.A2F_L_6_2(fpgaio_data_22_i),
.A2F_L_6_3(fpgaio_data_23_i),
.A2F_L_6_4(fpgaio_data_24_i),
.A2F_L_6_5(fpgaio_data_25_i),
.A2F_L_6_6(fpgaio_data_26_i),
.A2F_L_6_7(fpgaio_data_27_i),
.A2F_L_7_0(udma_cfg_data_30_i),
.A2F_L_7_1(udma_cfg_data_31_i),
.A2F_L_7_2(fpgaio_data_16_i),
.A2F_L_7_3(fpgaio_data_17_i),
.A2F_L_7_4(fpgaio_data_18_i),
.A2F_L_7_5(fpgaio_data_19_i),
.A2F_L_8_0(udma_cfg_data_22_i),
.A2F_L_8_1(udma_cfg_data_23_i),
.A2F_L_8_2(udma_cfg_data_24_i),
.A2F_L_8_3(udma_cfg_data_25_i),
.A2F_L_8_4(udma_cfg_data_26_i),
.A2F_L_8_5(udma_cfg_data_27_i),
.A2F_L_8_6(udma_cfg_data_28_i),
.A2F_L_8_7(udma_cfg_data_29_i),
.A2F_L_9_0(udma_cfg_data_16_i),
.A2F_L_9_1(udma_cfg_data_17_i),
.A2F_L_9_2(udma_cfg_data_18_i),
.A2F_L_9_3(udma_cfg_data_19_i),
.A2F_L_9_4(udma_cfg_data_20_i),
.A2F_L_9_5(udma_cfg_data_21_i),
.A2F_R_10_0(tcdm_r_rdata_p3_8_i),
.A2F_R_10_1(tcdm_r_rdata_p3_9_i),
.A2F_R_10_2(tcdm_r_rdata_p3_10_i),
.A2F_R_10_3(tcdm_r_rdata_p3_11_i),
.A2F_R_10_4(tcdm_r_rdata_p3_12_i),
.A2F_R_10_5(tcdm_r_rdata_p3_13_i),
.A2F_R_10_6(tcdm_r_rdata_p3_14_i),
.A2F_R_10_7(tcdm_r_rdata_p3_15_i),
.A2F_R_11_0(tcdm_r_rdata_p3_2_i),
.A2F_R_11_1(tcdm_r_rdata_p3_3_i),
.A2F_R_11_2(tcdm_r_rdata_p3_4_i),
.A2F_R_11_3(tcdm_r_rdata_p3_5_i),
.A2F_R_11_4(tcdm_r_rdata_p3_6_i),
.A2F_R_11_5(tcdm_r_rdata_p3_7_i),
.A2F_R_12_0(tcdm_r_rdata_p2_28_i),
.A2F_R_12_1(tcdm_r_rdata_p2_29_i),
.A2F_R_12_2(tcdm_r_rdata_p2_30_i),
.A2F_R_12_3(tcdm_r_rdata_p2_31_i),
.A2F_R_12_4(tcdm_gnt_p2_i),
.A2F_R_12_5(tcdm_r_valid_p2_i),
.A2F_R_12_6(tcdm_r_rdata_p3_0_i),
.A2F_R_12_7(tcdm_r_rdata_p3_1_i),
.A2F_R_13_0(tcdm_r_rdata_p2_22_i),
.A2F_R_13_1(tcdm_r_rdata_p2_23_i),
.A2F_R_13_2(tcdm_r_rdata_p2_24_i),
.A2F_R_13_3(tcdm_r_rdata_p2_25_i),
.A2F_R_13_4(tcdm_r_rdata_p2_26_i),
.A2F_R_13_5(tcdm_r_rdata_p2_27_i),
.A2F_R_14_0(tcdm_r_rdata_p2_14_i),
.A2F_R_14_1(tcdm_r_rdata_p2_15_i),
.A2F_R_14_2(tcdm_r_rdata_p2_16_i),
.A2F_R_14_3(tcdm_r_rdata_p2_17_i),
.A2F_R_14_4(tcdm_r_rdata_p2_18_i),
.A2F_R_14_5(tcdm_r_rdata_p2_19_i),
.A2F_R_14_6(tcdm_r_rdata_p2_20_i),
.A2F_R_14_7(tcdm_r_rdata_p2_21_i),
.A2F_R_15_0(tcdm_r_rdata_p2_8_i),
.A2F_R_15_1(tcdm_r_rdata_p2_9_i),
.A2F_R_15_2(tcdm_r_rdata_p2_10_i),
.A2F_R_15_3(tcdm_r_rdata_p2_11_i),
.A2F_R_15_4(tcdm_r_rdata_p2_12_i),
.A2F_R_15_5(tcdm_r_rdata_p2_13_i),
.A2F_R_16_0(tcdm_r_rdata_p2_0_i),
.A2F_R_16_1(tcdm_r_rdata_p2_1_i),
.A2F_R_16_2(tcdm_r_rdata_p2_2_i),
.A2F_R_16_3(tcdm_r_rdata_p2_3_i),
.A2F_R_16_4(tcdm_r_rdata_p2_4_i),
.A2F_R_16_5(tcdm_r_rdata_p2_5_i),
.A2F_R_16_6(tcdm_r_rdata_p2_6_i),
.A2F_R_16_7(tcdm_r_rdata_p2_7_i),
.A2F_R_17_0(tcdm_r_rdata_p0_0_i),
.A2F_R_17_1(tcdm_r_rdata_p0_1_i),
.A2F_R_17_2(tcdm_r_rdata_p0_2_i),
.A2F_R_17_3(tcdm_r_rdata_p0_3_i),
.A2F_R_17_4(tcdm_r_rdata_p0_4_i),
.A2F_R_17_5(tcdm_r_rdata_p0_5_i),
.A2F_R_18_0(tcdm_r_rdata_p0_6_i),
.A2F_R_18_1(tcdm_r_rdata_p0_7_i),
.A2F_R_18_2(tcdm_r_rdata_p0_8_i),
.A2F_R_18_3(tcdm_r_rdata_p0_9_i),
.A2F_R_18_4(tcdm_r_rdata_p0_10_i),
.A2F_R_18_5(tcdm_r_rdata_p0_11_i),
.A2F_R_18_6(tcdm_r_rdata_p0_12_i),
.A2F_R_18_7(tcdm_r_rdata_p0_13_i),
.A2F_R_19_0(tcdm_r_rdata_p0_14_i),
.A2F_R_19_1(tcdm_r_rdata_p0_15_i),
.A2F_R_19_2(tcdm_r_rdata_p0_16_i),
.A2F_R_19_3(tcdm_r_rdata_p0_17_i),
.A2F_R_19_4(tcdm_r_rdata_p0_18_i),
.A2F_R_19_5(tcdm_r_rdata_p0_19_i),
.A2F_R_1_0(supplyBus[302]),
.A2F_R_1_1(supplyBus[303]),
.A2F_R_1_2(supplyBus[304]),
.A2F_R_1_3(supplyBus[305]),
.A2F_R_1_4(supplyBus[306]),
.A2F_R_1_5(supplyBus[307]),
.A2F_R_20_0(tcdm_r_rdata_p0_20_i),
.A2F_R_20_1(tcdm_r_rdata_p0_21_i),
.A2F_R_20_2(tcdm_r_rdata_p0_22_i),
.A2F_R_20_3(tcdm_r_rdata_p0_23_i),
.A2F_R_20_4(tcdm_r_rdata_p0_24_i),
.A2F_R_20_5(tcdm_r_rdata_p0_25_i),
.A2F_R_20_6(tcdm_r_rdata_p0_26_i),
.A2F_R_20_7(tcdm_r_rdata_p0_27_i),
.A2F_R_21_0(tcdm_r_rdata_p0_28_i),
.A2F_R_21_1(tcdm_r_rdata_p0_29_i),
.A2F_R_21_2(tcdm_r_rdata_p0_30_i),
.A2F_R_21_3(tcdm_r_rdata_p0_31_i),
.A2F_R_21_4(tcdm_gnt_p0_i),
.A2F_R_21_5(tcdm_r_valid_p0_i),
.A2F_R_22_0(tcdm_r_rdata_p1_0_i),
.A2F_R_22_1(tcdm_r_rdata_p1_1_i),
.A2F_R_22_2(tcdm_r_rdata_p1_2_i),
.A2F_R_22_3(tcdm_r_rdata_p1_3_i),
.A2F_R_22_4(tcdm_r_rdata_p1_4_i),
.A2F_R_22_5(tcdm_r_rdata_p1_5_i),
.A2F_R_22_6(tcdm_r_rdata_p1_6_i),
.A2F_R_22_7(tcdm_r_rdata_p1_7_i),
.A2F_R_23_0(tcdm_r_rdata_p1_8_i),
.A2F_R_23_1(tcdm_r_rdata_p1_9_i),
.A2F_R_23_2(tcdm_r_rdata_p1_10_i),
.A2F_R_23_3(tcdm_r_rdata_p1_11_i),
.A2F_R_23_4(tcdm_r_rdata_p1_12_i),
.A2F_R_23_5(tcdm_r_rdata_p1_13_i),
.A2F_R_24_0(tcdm_r_rdata_p1_14_i),
.A2F_R_24_1(tcdm_r_rdata_p1_15_i),
.A2F_R_24_2(tcdm_r_rdata_p1_16_i),
.A2F_R_24_3(tcdm_r_rdata_p1_17_i),
.A2F_R_24_4(tcdm_r_rdata_p1_18_i),
.A2F_R_24_5(tcdm_r_rdata_p1_19_i),
.A2F_R_24_6(tcdm_r_rdata_p1_20_i),
.A2F_R_24_7(tcdm_r_rdata_p1_21_i),
.A2F_R_25_0(tcdm_r_rdata_p1_22_i),
.A2F_R_25_1(tcdm_r_rdata_p1_23_i),
.A2F_R_25_2(tcdm_r_rdata_p1_24_i),
.A2F_R_25_3(tcdm_r_rdata_p1_25_i),
.A2F_R_25_4(tcdm_r_rdata_p1_26_i),
.A2F_R_25_5(tcdm_r_rdata_p1_27_i),
.A2F_R_26_0(tcdm_r_rdata_p1_28_i),
.A2F_R_26_1(tcdm_r_rdata_p1_29_i),
.A2F_R_26_2(tcdm_r_rdata_p1_30_i),
.A2F_R_26_3(tcdm_r_rdata_p1_31_i),
.A2F_R_26_4(tcdm_gnt_p1_i),
.A2F_R_26_5(tcdm_r_valid_p1_i),
.A2F_R_26_6(fpgaio_data_8_i),
.A2F_R_26_7(fpgaio_data_9_i),
.A2F_R_27_0(fpgaio_data_10_i),
.A2F_R_27_1(fpgaio_data_11_i),
.A2F_R_27_2(RESET_RB),
.A2F_R_27_3(supplyBus[308]),
.A2F_R_27_4(supplyBus[309]),
.A2F_R_27_5(supplyBus[310]),
.A2F_R_28_0(supplyBus[311]),
.A2F_R_28_1(supplyBus[312]),
.A2F_R_28_2(supplyBus[313]),
.A2F_R_28_3(supplyBus[314]),
.A2F_R_28_4(supplyBus[315]),
.A2F_R_28_5(supplyBus[316]),
.A2F_R_28_6(supplyBus[317]),
.A2F_R_28_7(supplyBus[318]),
.A2F_R_29_0(supplyBus[319]),
.A2F_R_29_1(supplyBus[320]),
.A2F_R_29_2(supplyBus[321]),
.A2F_R_29_3(supplyBus[322]),
.A2F_R_29_4(supplyBus[323]),
.A2F_R_29_5(supplyBus[324]),
.A2F_R_2_0(supplyBus[325]),
.A2F_R_2_1(supplyBus[326]),
.A2F_R_2_2(supplyBus[327]),
.A2F_R_2_3(supplyBus[328]),
.A2F_R_2_4(supplyBus[329]),
.A2F_R_2_5(supplyBus[330]),
.A2F_R_2_6(supplyBus[331]),
.A2F_R_2_7(supplyBus[332]),
.A2F_R_30_0(supplyBus[333]),
.A2F_R_30_1(supplyBus[334]),
.A2F_R_30_2(supplyBus[335]),
.A2F_R_30_3(supplyBus[336]),
.A2F_R_30_4(supplyBus[337]),
.A2F_R_30_5(supplyBus[338]),
.A2F_R_30_6(supplyBus[339]),
.A2F_R_30_7(supplyBus[340]),
.A2F_R_31_0(supplyBus[341]),
.A2F_R_31_1(supplyBus[342]),
.A2F_R_31_2(supplyBus[343]),
.A2F_R_31_3(supplyBus[344]),
.A2F_R_31_4(supplyBus[345]),
.A2F_R_31_5(supplyBus[346]),
.A2F_R_32_0(supplyBus[347]),
.A2F_R_32_1(supplyBus[348]),
.A2F_R_32_2(supplyBus[349]),
.A2F_R_32_3(supplyBus[350]),
.A2F_R_32_4(supplyBus[351]),
.A2F_R_32_5(supplyBus[352]),
.A2F_R_32_6(supplyBus[353]),
.A2F_R_32_7(supplyBus[354]),
.A2F_R_3_0(supplyBus[355]),
.A2F_R_3_1(supplyBus[356]),
.A2F_R_3_2(supplyBus[357]),
.A2F_R_3_3(supplyBus[358]),
.A2F_R_3_4(supplyBus[359]),
.A2F_R_3_5(supplyBus[360]),
.A2F_R_4_0(supplyBus[361]),
.A2F_R_4_1(supplyBus[362]),
.A2F_R_4_2(supplyBus[363]),
.A2F_R_4_3(supplyBus[364]),
.A2F_R_4_4(supplyBus[365]),
.A2F_R_4_5(supplyBus[366]),
.A2F_R_4_6(supplyBus[367]),
.A2F_R_4_7(supplyBus[368]),
.A2F_R_5_0(supplyBus[369]),
.A2F_R_5_1(supplyBus[370]),
.A2F_R_5_2(supplyBus[371]),
.A2F_R_5_3(supplyBus[372]),
.A2F_R_5_4(supplyBus[373]),
.A2F_R_5_5(supplyBus[374]),
.A2F_R_6_0(fpgaio_data_14_i),
.A2F_R_6_1(fpgaio_data_15_i),
.A2F_R_6_2(RESET_RT),
.A2F_R_6_3(supplyBus[375]),
.A2F_R_6_4(supplyBus[376]),
.A2F_R_6_5(supplyBus[377]),
.A2F_R_6_6(supplyBus[378]),
.A2F_R_6_7(supplyBus[379]),
.A2F_R_7_0(tcdm_r_rdata_p3_30_i),
.A2F_R_7_1(tcdm_r_rdata_p3_31_i),
.A2F_R_7_2(tcdm_gnt_p3_i),
.A2F_R_7_3(tcdm_r_valid_p3_i),
.A2F_R_7_4(fpgaio_data_12_i),
.A2F_R_7_5(fpgaio_data_13_i),
.A2F_R_8_0(tcdm_r_rdata_p3_22_i),
.A2F_R_8_1(tcdm_r_rdata_p3_23_i),
.A2F_R_8_2(tcdm_r_rdata_p3_24_i),
.A2F_R_8_3(tcdm_r_rdata_p3_25_i),
.A2F_R_8_4(tcdm_r_rdata_p3_26_i),
.A2F_R_8_5(tcdm_r_rdata_p3_27_i),
.A2F_R_8_6(tcdm_r_rdata_p3_28_i),
.A2F_R_8_7(tcdm_r_rdata_p3_29_i),
.A2F_R_9_0(tcdm_r_rdata_p3_16_i),
.A2F_R_9_1(tcdm_r_rdata_p3_17_i),
.A2F_R_9_2(tcdm_r_rdata_p3_18_i),
.A2F_R_9_3(tcdm_r_rdata_p3_19_i),
.A2F_R_9_4(tcdm_r_rdata_p3_20_i),
.A2F_R_9_5(tcdm_r_rdata_p3_21_i),
.A2F_T_10_0(MU0_MATHB_EFPGA_MAC_OUT_7_),
.A2F_T_10_1(MU0_MATHB_EFPGA_MAC_OUT_6_),
.A2F_T_10_2(MU0_MATHB_EFPGA_MAC_OUT_5_),
.A2F_T_10_3(MU0_MATHB_EFPGA_MAC_OUT_4_),
.A2F_T_10_4(MU0_MATHB_EFPGA_MAC_OUT_3_),
.A2F_T_10_5(MU0_MATHB_EFPGA_MAC_OUT_2_),
.A2F_T_10_6(MU0_MATHB_EFPGA_MAC_OUT_1_),
.A2F_T_10_7(MU0_MATHB_EFPGA_MAC_OUT_0_),
.A2F_T_11_0(supplyBus[380]),
.A2F_T_11_1(supplyBus[381]),
.A2F_T_11_2(MU0_TPRAM_EFPGA_COEF_R_DATA_31_),
.A2F_T_11_3(MU0_TPRAM_EFPGA_COEF_R_DATA_30_),
.A2F_T_11_4(MU0_TPRAM_EFPGA_COEF_R_DATA_29_),
.A2F_T_11_5(MU0_TPRAM_EFPGA_COEF_R_DATA_28_),
.A2F_T_12_0(MU0_TPRAM_EFPGA_COEF_R_DATA_27_),
.A2F_T_12_1(MU0_TPRAM_EFPGA_COEF_R_DATA_26_),
.A2F_T_12_2(MU0_TPRAM_EFPGA_COEF_R_DATA_25_),
.A2F_T_12_3(MU0_TPRAM_EFPGA_COEF_R_DATA_24_),
.A2F_T_12_4(MU0_TPRAM_EFPGA_COEF_R_DATA_23_),
.A2F_T_12_5(MU0_TPRAM_EFPGA_COEF_R_DATA_22_),
.A2F_T_12_6(MU0_TPRAM_EFPGA_COEF_R_DATA_21_),
.A2F_T_12_7(MU0_TPRAM_EFPGA_COEF_R_DATA_20_),
.A2F_T_13_0(MU0_TPRAM_EFPGA_COEF_R_DATA_19_),
.A2F_T_13_1(MU0_TPRAM_EFPGA_COEF_R_DATA_18_),
.A2F_T_13_2(MU0_TPRAM_EFPGA_COEF_R_DATA_17_),
.A2F_T_13_3(MU0_TPRAM_EFPGA_COEF_R_DATA_16_),
.A2F_T_13_4(MU0_TPRAM_EFPGA_COEF_R_DATA_15_),
.A2F_T_13_5(MU0_TPRAM_EFPGA_COEF_R_DATA_14_),
.A2F_T_14_0(MU0_TPRAM_EFPGA_COEF_R_DATA_13_),
.A2F_T_14_1(MU0_TPRAM_EFPGA_COEF_R_DATA_12_),
.A2F_T_14_2(MU0_TPRAM_EFPGA_COEF_R_DATA_11_),
.A2F_T_14_3(MU0_TPRAM_EFPGA_COEF_R_DATA_10_),
.A2F_T_14_4(MU0_TPRAM_EFPGA_COEF_R_DATA_9_),
.A2F_T_14_5(MU0_TPRAM_EFPGA_COEF_R_DATA_8_),
.A2F_T_14_6(MU0_TPRAM_EFPGA_COEF_R_DATA_7_),
.A2F_T_14_7(MU0_TPRAM_EFPGA_COEF_R_DATA_6_),
.A2F_T_15_0(MU0_TPRAM_EFPGA_COEF_R_DATA_5_),
.A2F_T_15_1(MU0_TPRAM_EFPGA_COEF_R_DATA_4_),
.A2F_T_15_2(MU0_TPRAM_EFPGA_COEF_R_DATA_3_),
.A2F_T_15_3(MU0_TPRAM_EFPGA_COEF_R_DATA_2_),
.A2F_T_15_4(MU0_TPRAM_EFPGA_COEF_R_DATA_1_),
.A2F_T_15_5(MU0_TPRAM_EFPGA_COEF_R_DATA_0_),
.A2F_T_16_0(supplyBus[382]),
.A2F_T_16_1(supplyBus[383]),
.A2F_T_16_2(supplyBus[384]),
.A2F_T_16_3(supplyBus[385]),
.A2F_T_16_4(supplyBus[386]),
.A2F_T_16_5(supplyBus[387]),
.A2F_T_16_6(supplyBus[388]),
.A2F_T_16_7(supplyBus[389]),
.A2F_T_17_0(MU1_TPRAM_EFPGA_OPER_R_DATA_31_),
.A2F_T_17_1(MU1_TPRAM_EFPGA_OPER_R_DATA_30_),
.A2F_T_17_2(MU1_TPRAM_EFPGA_OPER_R_DATA_29_),
.A2F_T_17_3(MU1_TPRAM_EFPGA_OPER_R_DATA_28_),
.A2F_T_17_4(MU1_TPRAM_EFPGA_OPER_R_DATA_27_),
.A2F_T_17_5(MU1_TPRAM_EFPGA_OPER_R_DATA_26_),
.A2F_T_18_0(MU1_TPRAM_EFPGA_OPER_R_DATA_25_),
.A2F_T_18_1(MU1_TPRAM_EFPGA_OPER_R_DATA_24_),
.A2F_T_18_2(MU1_TPRAM_EFPGA_OPER_R_DATA_23_),
.A2F_T_18_3(MU1_TPRAM_EFPGA_OPER_R_DATA_22_),
.A2F_T_18_4(MU1_TPRAM_EFPGA_OPER_R_DATA_21_),
.A2F_T_18_5(MU1_TPRAM_EFPGA_OPER_R_DATA_20_),
.A2F_T_18_6(MU1_TPRAM_EFPGA_OPER_R_DATA_19_),
.A2F_T_18_7(MU1_TPRAM_EFPGA_OPER_R_DATA_18_),
.A2F_T_19_0(MU1_TPRAM_EFPGA_OPER_R_DATA_17_),
.A2F_T_19_1(MU1_TPRAM_EFPGA_OPER_R_DATA_16_),
.A2F_T_19_2(MU1_TPRAM_EFPGA_OPER_R_DATA_15_),
.A2F_T_19_3(MU1_TPRAM_EFPGA_OPER_R_DATA_14_),
.A2F_T_19_4(MU1_TPRAM_EFPGA_OPER_R_DATA_13_),
.A2F_T_19_5(MU1_TPRAM_EFPGA_OPER_R_DATA_12_),
.A2F_T_1_0(supplyBus[390]),
.A2F_T_1_1(supplyBus[391]),
.A2F_T_1_2(MU0_TPRAM_EFPGA_OPER_R_DATA_31_),
.A2F_T_1_3(MU0_TPRAM_EFPGA_OPER_R_DATA_30_),
.A2F_T_1_4(MU0_TPRAM_EFPGA_OPER_R_DATA_29_),
.A2F_T_1_5(MU0_TPRAM_EFPGA_OPER_R_DATA_28_),
.A2F_T_20_0(MU1_TPRAM_EFPGA_OPER_R_DATA_11_),
.A2F_T_20_1(MU1_TPRAM_EFPGA_OPER_R_DATA_10_),
.A2F_T_20_2(MU1_TPRAM_EFPGA_OPER_R_DATA_9_),
.A2F_T_20_3(MU1_TPRAM_EFPGA_OPER_R_DATA_8_),
.A2F_T_20_4(MU1_TPRAM_EFPGA_OPER_R_DATA_7_),
.A2F_T_20_5(MU1_TPRAM_EFPGA_OPER_R_DATA_6_),
.A2F_T_20_6(MU1_TPRAM_EFPGA_OPER_R_DATA_5_),
.A2F_T_20_7(MU1_TPRAM_EFPGA_OPER_R_DATA_4_),
.A2F_T_21_0(MU1_TPRAM_EFPGA_OPER_R_DATA_3_),
.A2F_T_21_1(MU1_TPRAM_EFPGA_OPER_R_DATA_2_),
.A2F_T_21_2(MU1_TPRAM_EFPGA_OPER_R_DATA_1_),
.A2F_T_21_3(MU1_TPRAM_EFPGA_OPER_R_DATA_0_),
.A2F_T_21_4(supplyBus[392]),
.A2F_T_21_5(supplyBus[393]),
.A2F_T_22_0(supplyBus[394]),
.A2F_T_22_1(supplyBus[395]),
.A2F_T_22_2(supplyBus[396]),
.A2F_T_22_3(supplyBus[397]),
.A2F_T_22_4(supplyBus[398]),
.A2F_T_22_5(supplyBus[399]),
.A2F_T_22_6(supplyBus[400]),
.A2F_T_22_7(supplyBus[401]),
.A2F_T_23_0(MU1_MATHB_EFPGA_MAC_OUT_31_),
.A2F_T_23_1(MU1_MATHB_EFPGA_MAC_OUT_30_),
.A2F_T_23_2(MU1_MATHB_EFPGA_MAC_OUT_29_),
.A2F_T_23_3(MU1_MATHB_EFPGA_MAC_OUT_28_),
.A2F_T_23_4(MU1_MATHB_EFPGA_MAC_OUT_27_),
.A2F_T_23_5(MU1_MATHB_EFPGA_MAC_OUT_26_),
.A2F_T_24_0(MU1_MATHB_EFPGA_MAC_OUT_25_),
.A2F_T_24_1(MU1_MATHB_EFPGA_MAC_OUT_24_),
.A2F_T_24_2(MU1_MATHB_EFPGA_MAC_OUT_23_),
.A2F_T_24_3(MU1_MATHB_EFPGA_MAC_OUT_22_),
.A2F_T_24_4(MU1_MATHB_EFPGA_MAC_OUT_21_),
.A2F_T_24_5(MU1_MATHB_EFPGA_MAC_OUT_20_),
.A2F_T_24_6(MU1_MATHB_EFPGA_MAC_OUT_19_),
.A2F_T_24_7(MU1_MATHB_EFPGA_MAC_OUT_18_),
.A2F_T_25_0(MU1_MATHB_EFPGA_MAC_OUT_17_),
.A2F_T_25_1(MU1_MATHB_EFPGA_MAC_OUT_16_),
.A2F_T_25_2(MU1_MATHB_EFPGA_MAC_OUT_15_),
.A2F_T_25_3(MU1_MATHB_EFPGA_MAC_OUT_14_),
.A2F_T_25_4(MU1_MATHB_EFPGA_MAC_OUT_13_),
.A2F_T_25_5(MU1_MATHB_EFPGA_MAC_OUT_12_),
.A2F_T_26_0(MU1_MATHB_EFPGA_MAC_OUT_11_),
.A2F_T_26_1(MU1_MATHB_EFPGA_MAC_OUT_10_),
.A2F_T_26_2(MU1_MATHB_EFPGA_MAC_OUT_9_),
.A2F_T_26_3(MU1_MATHB_EFPGA_MAC_OUT_8_),
.A2F_T_26_4(MU1_MATHB_EFPGA_MAC_OUT_7_),
.A2F_T_26_5(MU1_MATHB_EFPGA_MAC_OUT_6_),
.A2F_T_26_6(MU1_MATHB_EFPGA_MAC_OUT_5_),
.A2F_T_26_7(MU1_MATHB_EFPGA_MAC_OUT_4_),
.A2F_T_27_0(MU1_MATHB_EFPGA_MAC_OUT_3_),
.A2F_T_27_1(MU1_MATHB_EFPGA_MAC_OUT_2_),
.A2F_T_27_2(MU1_MATHB_EFPGA_MAC_OUT_1_),
.A2F_T_27_3(MU1_MATHB_EFPGA_MAC_OUT_0_),
.A2F_T_27_4(supplyBus[402]),
.A2F_T_27_5(supplyBus[403]),
.A2F_T_28_0(MU1_TPRAM_EFPGA_COEF_R_DATA_31_),
.A2F_T_28_1(MU1_TPRAM_EFPGA_COEF_R_DATA_30_),
.A2F_T_28_2(MU1_TPRAM_EFPGA_COEF_R_DATA_29_),
.A2F_T_28_3(MU1_TPRAM_EFPGA_COEF_R_DATA_28_),
.A2F_T_28_4(MU1_TPRAM_EFPGA_COEF_R_DATA_27_),
.A2F_T_28_5(MU1_TPRAM_EFPGA_COEF_R_DATA_26_),
.A2F_T_28_6(MU1_TPRAM_EFPGA_COEF_R_DATA_25_),
.A2F_T_28_7(MU1_TPRAM_EFPGA_COEF_R_DATA_24_),
.A2F_T_29_0(MU1_TPRAM_EFPGA_COEF_R_DATA_23_),
.A2F_T_29_1(MU1_TPRAM_EFPGA_COEF_R_DATA_22_),
.A2F_T_29_2(MU1_TPRAM_EFPGA_COEF_R_DATA_21_),
.A2F_T_29_3(MU1_TPRAM_EFPGA_COEF_R_DATA_20_),
.A2F_T_29_4(MU1_TPRAM_EFPGA_COEF_R_DATA_19_),
.A2F_T_29_5(MU1_TPRAM_EFPGA_COEF_R_DATA_18_),
.A2F_T_2_0(MU0_TPRAM_EFPGA_OPER_R_DATA_27_),
.A2F_T_2_1(MU0_TPRAM_EFPGA_OPER_R_DATA_26_),
.A2F_T_2_2(MU0_TPRAM_EFPGA_OPER_R_DATA_25_),
.A2F_T_2_3(MU0_TPRAM_EFPGA_OPER_R_DATA_24_),
.A2F_T_2_4(MU0_TPRAM_EFPGA_OPER_R_DATA_23_),
.A2F_T_2_5(MU0_TPRAM_EFPGA_OPER_R_DATA_22_),
.A2F_T_2_6(MU0_TPRAM_EFPGA_OPER_R_DATA_21_),
.A2F_T_2_7(MU0_TPRAM_EFPGA_OPER_R_DATA_20_),
.A2F_T_30_0(MU1_TPRAM_EFPGA_COEF_R_DATA_17_),
.A2F_T_30_1(MU1_TPRAM_EFPGA_COEF_R_DATA_16_),
.A2F_T_30_2(MU1_TPRAM_EFPGA_COEF_R_DATA_15_),
.A2F_T_30_3(MU1_TPRAM_EFPGA_COEF_R_DATA_14_),
.A2F_T_30_4(MU1_TPRAM_EFPGA_COEF_R_DATA_13_),
.A2F_T_30_5(MU1_TPRAM_EFPGA_COEF_R_DATA_12_),
.A2F_T_30_6(MU1_TPRAM_EFPGA_COEF_R_DATA_11_),
.A2F_T_30_7(MU1_TPRAM_EFPGA_COEF_R_DATA_10_),
.A2F_T_31_0(MU1_TPRAM_EFPGA_COEF_R_DATA_9_),
.A2F_T_31_1(MU1_TPRAM_EFPGA_COEF_R_DATA_8_),
.A2F_T_31_2(MU1_TPRAM_EFPGA_COEF_R_DATA_7_),
.A2F_T_31_3(MU1_TPRAM_EFPGA_COEF_R_DATA_6_),
.A2F_T_31_4(MU1_TPRAM_EFPGA_COEF_R_DATA_5_),
.A2F_T_31_5(MU1_TPRAM_EFPGA_COEF_R_DATA_4_),
.A2F_T_32_0(MU1_TPRAM_EFPGA_COEF_R_DATA_3_),
.A2F_T_32_1(MU1_TPRAM_EFPGA_COEF_R_DATA_2_),
.A2F_T_32_2(MU1_TPRAM_EFPGA_COEF_R_DATA_1_),
.A2F_T_32_3(MU1_TPRAM_EFPGA_COEF_R_DATA_0_),
.A2F_T_32_4(supplyBus[404]),
.A2F_T_32_5(supplyBus[405]),
.A2F_T_32_6(supplyBus[406]),
.A2F_T_32_7(supplyBus[407]),
.A2F_T_3_0(MU0_TPRAM_EFPGA_OPER_R_DATA_19_),
.A2F_T_3_1(MU0_TPRAM_EFPGA_OPER_R_DATA_18_),
.A2F_T_3_2(MU0_TPRAM_EFPGA_OPER_R_DATA_17_),
.A2F_T_3_3(MU0_TPRAM_EFPGA_OPER_R_DATA_16_),
.A2F_T_3_4(MU0_TPRAM_EFPGA_OPER_R_DATA_15_),
.A2F_T_3_5(MU0_TPRAM_EFPGA_OPER_R_DATA_14_),
.A2F_T_4_0(MU0_TPRAM_EFPGA_OPER_R_DATA_13_),
.A2F_T_4_1(MU0_TPRAM_EFPGA_OPER_R_DATA_12_),
.A2F_T_4_2(MU0_TPRAM_EFPGA_OPER_R_DATA_11_),
.A2F_T_4_3(MU0_TPRAM_EFPGA_OPER_R_DATA_10_),
.A2F_T_4_4(MU0_TPRAM_EFPGA_OPER_R_DATA_9_),
.A2F_T_4_5(MU0_TPRAM_EFPGA_OPER_R_DATA_8_),
.A2F_T_4_6(MU0_TPRAM_EFPGA_OPER_R_DATA_7_),
.A2F_T_4_7(MU0_TPRAM_EFPGA_OPER_R_DATA_6_),
.A2F_T_5_0(MU0_TPRAM_EFPGA_OPER_R_DATA_5_),
.A2F_T_5_1(MU0_TPRAM_EFPGA_OPER_R_DATA_4_),
.A2F_T_5_2(MU0_TPRAM_EFPGA_OPER_R_DATA_3_),
.A2F_T_5_3(MU0_TPRAM_EFPGA_OPER_R_DATA_2_),
.A2F_T_5_4(MU0_TPRAM_EFPGA_OPER_R_DATA_1_),
.A2F_T_5_5(MU0_TPRAM_EFPGA_OPER_R_DATA_0_),
.A2F_T_6_0(supplyBus[408]),
.A2F_T_6_1(supplyBus[409]),
.A2F_T_6_2(supplyBus[410]),
.A2F_T_6_3(supplyBus[411]),
.A2F_T_6_4(MU0_MATHB_EFPGA_MAC_OUT_31_),
.A2F_T_6_5(MU0_MATHB_EFPGA_MAC_OUT_30_),
.A2F_T_6_6(MU0_MATHB_EFPGA_MAC_OUT_29_),
.A2F_T_6_7(MU0_MATHB_EFPGA_MAC_OUT_28_),
.A2F_T_7_0(MU0_MATHB_EFPGA_MAC_OUT_27_),
.A2F_T_7_1(MU0_MATHB_EFPGA_MAC_OUT_26_),
.A2F_T_7_2(MU0_MATHB_EFPGA_MAC_OUT_25_),
.A2F_T_7_3(MU0_MATHB_EFPGA_MAC_OUT_24_),
.A2F_T_7_4(MU0_MATHB_EFPGA_MAC_OUT_23_),
.A2F_T_7_5(MU0_MATHB_EFPGA_MAC_OUT_22_),
.A2F_T_8_0(MU0_MATHB_EFPGA_MAC_OUT_21_),
.A2F_T_8_1(MU0_MATHB_EFPGA_MAC_OUT_20_),
.A2F_T_8_2(MU0_MATHB_EFPGA_MAC_OUT_19_),
.A2F_T_8_3(MU0_MATHB_EFPGA_MAC_OUT_18_),
.A2F_T_8_4(MU0_MATHB_EFPGA_MAC_OUT_17_),
.A2F_T_8_5(MU0_MATHB_EFPGA_MAC_OUT_16_),
.A2F_T_8_6(MU0_MATHB_EFPGA_MAC_OUT_15_),
.A2F_T_8_7(MU0_MATHB_EFPGA_MAC_OUT_14_),
.A2F_T_9_0(MU0_MATHB_EFPGA_MAC_OUT_13_),
.A2F_T_9_1(MU0_MATHB_EFPGA_MAC_OUT_12_),
.A2F_T_9_2(MU0_MATHB_EFPGA_MAC_OUT_11_),
.A2F_T_9_3(MU0_MATHB_EFPGA_MAC_OUT_10_),
.A2F_T_9_4(MU0_MATHB_EFPGA_MAC_OUT_9_),
.A2F_T_9_5(MU0_MATHB_EFPGA_MAC_OUT_8_),
.A2Freg_B_11_0(supplyBus[412]),
.A2Freg_B_13_0(supplyBus[413]),
.A2Freg_B_15_0(supplyBus[414]),
.A2Freg_B_17_0(supplyBus[415]),
.A2Freg_B_19_0(supplyBus[416]),
.A2Freg_B_1_0(supplyBus[417]),
.A2Freg_B_21_0(supplyBus[418]),
.A2Freg_B_23_0(supplyBus[419]),
.A2Freg_B_25_0(supplyBus[420]),
.A2Freg_B_27_0(supplyBus[421]),
.A2Freg_B_29_0(supplyBus[422]),
.A2Freg_B_31_0(supplyBus[423]),
.A2Freg_B_3_0(supplyBus[424]),
.A2Freg_B_5_0(supplyBus[425]),
.A2Freg_B_7_0(supplyBus[426]),
.A2Freg_B_9_0(supplyBus[427]),
.A2Freg_L_11_0(supplyBus[428]),
.A2Freg_L_13_0(supplyBus[429]),
.A2Freg_L_15_0(supplyBus[430]),
.A2Freg_L_17_0(supplyBus[431]),
.A2Freg_L_19_0(supplyBus[432]),
.A2Freg_L_1_0(supplyBus[433]),
.A2Freg_L_21_0(supplyBus[434]),
.A2Freg_L_23_0(supplyBus[435]),
.A2Freg_L_25_0(supplyBus[436]),
.A2Freg_L_27_0(supplyBus[437]),
.A2Freg_L_29_0(supplyBus[438]),
.A2Freg_L_31_0(supplyBus[439]),
.A2Freg_L_3_0(supplyBus[440]),
.A2Freg_L_5_0(supplyBus[441]),
.A2Freg_L_7_0(supplyBus[442]),
.A2Freg_L_9_0(supplyBus[443]),
.A2Freg_R_11_0(supplyBus[444]),
.A2Freg_R_13_0(supplyBus[445]),
.A2Freg_R_15_0(supplyBus[446]),
.A2Freg_R_17_0(supplyBus[447]),
.A2Freg_R_19_0(supplyBus[448]),
.A2Freg_R_1_0(supplyBus[449]),
.A2Freg_R_21_0(supplyBus[450]),
.A2Freg_R_23_0(supplyBus[451]),
.A2Freg_R_25_0(supplyBus[452]),
.A2Freg_R_27_0(supplyBus[453]),
.A2Freg_R_29_0(supplyBus[454]),
.A2Freg_R_31_0(supplyBus[455]),
.A2Freg_R_3_0(supplyBus[456]),
.A2Freg_R_5_0(supplyBus[457]),
.A2Freg_R_7_0(supplyBus[458]),
.A2Freg_R_9_0(supplyBus[459]),
.A2Freg_T_11_0(supplyBus[460]),
.A2Freg_T_13_0(supplyBus[461]),
.A2Freg_T_15_0(supplyBus[462]),
.A2Freg_T_17_0(supplyBus[463]),
.A2Freg_T_19_0(supplyBus[464]),
.A2Freg_T_1_0(supplyBus[465]),
.A2Freg_T_21_0(supplyBus[466]),
.A2Freg_T_23_0(supplyBus[467]),
.A2Freg_T_25_0(supplyBus[468]),
.A2Freg_T_27_0(supplyBus[469]),
.A2Freg_T_29_0(supplyBus[470]),
.A2Freg_T_31_0(supplyBus[471]),
.A2Freg_T_3_0(supplyBus[472]),
.A2Freg_T_5_0(supplyBus[473]),
.A2Freg_T_7_0(supplyBus[474]),
.A2Freg_T_9_0(supplyBus[475]),
. M_0_( M_0_),
.BL_CLK(BL_CLK),
.BL_DIN_0_(BL_DIN_0_),
.BL_DIN_10_(BL_DIN_10_),
.BL_DIN_11_(BL_DIN_11_),
.BL_DIN_12_(BL_DIN_12_),
.BL_DIN_13_(BL_DIN_13_),
.BL_DIN_14_(BL_DIN_14_),
.BL_DIN_15_(BL_DIN_15_),
.BL_DIN_16_(BL_DIN_16_),
.BL_DIN_17_(BL_DIN_17_),
.BL_DIN_18_(BL_DIN_18_),
.BL_DIN_19_(BL_DIN_19_),
.BL_DIN_1_(BL_DIN_1_),
.BL_DIN_20_(BL_DIN_20_),
.BL_DIN_21_(BL_DIN_21_),
.BL_DIN_22_(BL_DIN_22_),
.BL_DIN_23_(BL_DIN_23_),
.BL_DIN_24_(BL_DIN_24_),
.BL_DIN_25_(BL_DIN_25_),
.BL_DIN_26_(BL_DIN_26_),
.BL_DIN_27_(BL_DIN_27_),
.BL_DIN_28_(BL_DIN_28_),
.BL_DIN_29_(BL_DIN_29_),
.BL_DIN_2_(BL_DIN_2_),
.BL_DIN_30_(BL_DIN_30_),
.BL_DIN_31_(BL_DIN_31_),
.BL_DIN_3_(BL_DIN_3_),
.BL_DIN_4_(BL_DIN_4_),
.BL_DIN_5_(BL_DIN_5_),
.BL_DIN_6_(BL_DIN_6_),
.BL_DIN_7_(BL_DIN_7_),
.BL_DIN_8_(BL_DIN_8_),
.BL_DIN_9_(BL_DIN_9_),
.BL_PWRGATE_0_(BL_PWRGATE_0_),
.BL_PWRGATE_1_(BL_PWRGATE_1_),
.BL_PWRGATE_2_(BL_PWRGATE_2_),
.BL_PWRGATE_3_(BL_PWRGATE_3_),
.CLOAD_DIN_SEL(CLOAD_DIN_SEL),
.DIN_INT_L_ONLY(DIN_INT_L_ONLY),
.DIN_INT_R_ONLY(DIN_INT_R_ONLY),
.DIN_SLC_TB_INT(DIN_SLC_TB_INT),
.FB_CFG_DONE(FB_CFG_DONE),
.FB_ISO_ENB(FB_ISO_ENB),
.FB_SPE_IN_0_(FB_SPE_IN_0_),
.FB_SPE_IN_1_(FB_SPE_IN_1_),
.FB_SPE_IN_2_(FB_SPE_IN_2_),
.FB_SPE_IN_3_(FB_SPE_IN_3_),
.ISO_EN_0_(ISO_EN_0_),
.ISO_EN_1_(ISO_EN_1_),
.ISO_EN_2_(ISO_EN_2_),
.ISO_EN_3_(ISO_EN_3_),
.MLATCH(MLATCH),
.M_1_(M_1_),
.M_2_(M_2_),
.M_3_(M_3_),
.M_4_(M_4_),
.M_5_(M_5_),
.NB(NB),
.PB(PB),
.PCHG_B(PCHG_B),
.PI_PWR_0_(PI_PWR_0_),
.PI_PWR_1_(PI_PWR_1_),
.PI_PWR_2_(PI_PWR_2_),
.PI_PWR_3_(PI_PWR_3_),
.POR(POR),
.PROG_0_(PROG_0_),
.PROG_1_(PROG_1_),
.PROG_2_(PROG_2_),
.PROG_3_(PROG_3_),
.PROG_IFX(PROG_IFX),
.PWR_GATE(PWR_GATE),
.RE(RE),
.STM(STM),
.VLP_CLKDIS_0_(VLP_CLKDIS_0_),
.VLP_CLKDIS_1_(VLP_CLKDIS_1_),
.VLP_CLKDIS_2_(VLP_CLKDIS_2_),
.VLP_CLKDIS_3_(VLP_CLKDIS_3_),
.VLP_CLKDIS_IFX(VLP_CLKDIS_IFX),
.VLP_PWRDIS_0_(VLP_PWRDIS_0_),
.VLP_PWRDIS_1_(VLP_PWRDIS_1_),
.VLP_PWRDIS_2_(VLP_PWRDIS_2_),
.VLP_PWRDIS_3_(VLP_PWRDIS_3_),
.VLP_PWRDIS_IFX(VLP_PWRDIS_IFX),
.VLP_SRDIS_0_(VLP_SRDIS_0_),
.VLP_SRDIS_1_(VLP_SRDIS_1_),
.VLP_SRDIS_2_(VLP_SRDIS_2_),
.VLP_SRDIS_3_(VLP_SRDIS_3_),
.VLP_SRDIS_IFX(VLP_SRDIS_IFX),
.WE(WE),
.WE_INT(WE_INT),
.WL_CLK(WL_CLK),
.WL_CLOAD_SEL_0_(WL_CLOAD_SEL_0_),
.WL_CLOAD_SEL_1_(WL_CLOAD_SEL_1_),
.WL_CLOAD_SEL_2_(WL_CLOAD_SEL_2_),
.WL_DIN_0_(WL_DIN_0_),
.WL_DIN_1_(WL_DIN_1_),
.WL_DIN_2_(WL_DIN_2_),
.WL_DIN_3_(WL_DIN_3_),
.WL_DIN_4_(WL_DIN_4_),
.WL_DIN_5_(WL_DIN_5_),
.WL_EN(WL_EN),
.WL_INT_DIN_SEL(WL_INT_DIN_SEL),
.WL_PWRGATE_0_(WL_PWRGATE_0_),
.WL_PWRGATE_1_(WL_PWRGATE_1_),
.WL_RESETB(WL_RESETB),
.WL_SEL_0_(WL_SEL_0_),
.WL_SEL_1_(WL_SEL_1_),
.WL_SEL_2_(WL_SEL_2_),
.WL_SEL_3_(WL_SEL_3_),
.WL_SEL_TB_INT(WL_SEL_TB_INT),
.F2A_B_10_0(),
.F2A_B_10_1(),
.F2A_B_10_10(),
.F2A_B_10_11(),
.F2A_B_10_12(),
.F2A_B_10_13(),
.F2A_B_10_14(),
.F2A_B_10_15(),
.F2A_B_10_16(),
.F2A_B_10_17(),
.F2A_B_10_2(),
.F2A_B_10_3(),
.F2A_B_10_4(),
.F2A_B_10_5(),
.F2A_B_10_6(),
.F2A_B_10_7(),
.F2A_B_10_8(),
.F2A_B_10_9(),
.F2A_B_11_0(),
.F2A_B_11_1(),
.F2A_B_11_10(),
.F2A_B_11_11(),
.F2A_B_11_2(),
.F2A_B_11_3(),
.F2A_B_11_4(),
.F2A_B_11_5(),
.F2A_B_11_6(),
.F2A_B_11_7(),
.F2A_B_11_8(),
.F2A_B_11_9(),
.F2A_B_12_0(),
.F2A_B_12_1(),
.F2A_B_12_10(),
.F2A_B_12_11(),
.F2A_B_12_12(),
.F2A_B_12_13(),
.F2A_B_12_14(),
.F2A_B_12_15(),
.F2A_B_12_16(),
.F2A_B_12_17(),
.F2A_B_12_2(),
.F2A_B_12_3(),
.F2A_B_12_4(),
.F2A_B_12_5(),
.F2A_B_12_6(),
.F2A_B_12_7(),
.F2A_B_12_8(),
.F2A_B_12_9(),
.F2A_B_13_0(),
.F2A_B_13_1(),
.F2A_B_13_10(),
.F2A_B_13_11(),
.F2A_B_13_2(),
.F2A_B_13_3(),
.F2A_B_13_4(),
.F2A_B_13_5(),
.F2A_B_13_6(),
.F2A_B_13_7(),
.F2A_B_13_8(),
.F2A_B_13_9(),
.F2A_B_14_0(),
.F2A_B_14_1(),
.F2A_B_14_10(),
.F2A_B_14_11(),
.F2A_B_14_12(),
.F2A_B_14_13(),
.F2A_B_14_14(),
.F2A_B_14_15(),
.F2A_B_14_16(),
.F2A_B_14_17(),
.F2A_B_14_2(),
.F2A_B_14_3(),
.F2A_B_14_4(),
.F2A_B_14_5(),
.F2A_B_14_6(),
.F2A_B_14_7(),
.F2A_B_14_8(),
.F2A_B_14_9(),
.F2A_B_15_0(),
.F2A_B_15_1(),
.F2A_B_15_10(),
.F2A_B_15_11(),
.F2A_B_15_2(),
.F2A_B_15_3(),
.F2A_B_15_4(),
.F2A_B_15_5(),
.F2A_B_15_6(),
.F2A_B_15_7(),
.F2A_B_15_8(),
.F2A_B_15_9(),
.F2A_B_16_0(fpgaio_oe_0_o),
.F2A_B_16_1(fpgaio_data_0_o),
.F2A_B_16_10(),
.F2A_B_16_11(),
.F2A_B_16_12(),
.F2A_B_16_13(),
.F2A_B_16_17(),
.F2A_B_16_2(fpgaio_oe_1_o),
.F2A_B_16_3(fpgaio_data_1_o),
.F2A_B_16_4(fpgaio_oe_2_o),
.F2A_B_16_5(fpgaio_data_2_o),
.F2A_B_16_6(fpgaio_oe_3_o),
.F2A_B_16_7(fpgaio_data_3_o),
.F2A_B_16_8(),
.F2A_B_16_9(),
.F2A_B_17_0(fpgaio_oe_4_o),
.F2A_B_17_1(fpgaio_data_4_o),
.F2A_B_17_10(),
.F2A_B_17_11(),
.F2A_B_17_2(fpgaio_oe_5_o),
.F2A_B_17_3(fpgaio_data_5_o),
.F2A_B_17_4(fpgaio_oe_6_o),
.F2A_B_17_5(fpgaio_data_6_o),
.F2A_B_17_6(fpgaio_oe_7_o),
.F2A_B_17_7(fpgaio_data_7_o),
.F2A_B_17_8(),
.F2A_B_17_9(),
.F2A_B_18_0(),
.F2A_B_18_1(),
.F2A_B_18_10(),
.F2A_B_18_11(),
.F2A_B_18_12(),
.F2A_B_18_13(),
.F2A_B_18_14(),
.F2A_B_18_15(),
.F2A_B_18_16(),
.F2A_B_18_17(),
.F2A_B_18_2(),
.F2A_B_18_3(),
.F2A_B_18_4(),
.F2A_B_18_5(),
.F2A_B_18_6(),
.F2A_B_18_7(),
.F2A_B_18_8(),
.F2A_B_18_9(),
.F2A_B_19_0(),
.F2A_B_19_1(),
.F2A_B_19_10(),
.F2A_B_19_11(),
.F2A_B_19_2(),
.F2A_B_19_3(),
.F2A_B_19_4(),
.F2A_B_19_5(),
.F2A_B_19_6(),
.F2A_B_19_7(),
.F2A_B_19_8(),
.F2A_B_19_9(),
.F2A_B_1_0(),
.F2A_B_1_1(),
.F2A_B_1_10(),
.F2A_B_1_11(),
.F2A_B_1_2(),
.F2A_B_1_3(),
.F2A_B_1_4(),
.F2A_B_1_5(),
.F2A_B_1_6(),
.F2A_B_1_7(),
.F2A_B_1_8(),
.F2A_B_1_9(),
.F2A_B_20_0(),
.F2A_B_20_1(),
.F2A_B_20_10(),
.F2A_B_20_11(),
.F2A_B_20_12(),
.F2A_B_20_13(),
.F2A_B_20_14(),
.F2A_B_20_15(),
.F2A_B_20_16(),
.F2A_B_20_17(),
.F2A_B_20_2(),
.F2A_B_20_3(),
.F2A_B_20_4(),
.F2A_B_20_5(),
.F2A_B_20_6(),
.F2A_B_20_7(),
.F2A_B_20_8(),
.F2A_B_20_9(),
.F2A_B_21_0(),
.F2A_B_21_1(),
.F2A_B_21_10(),
.F2A_B_21_11(),
.F2A_B_21_2(),
.F2A_B_21_3(),
.F2A_B_21_4(),
.F2A_B_21_5(),
.F2A_B_21_6(),
.F2A_B_21_7(),
.F2A_B_21_8(),
.F2A_B_21_9(),
.F2A_B_22_0(),
.F2A_B_22_1(),
.F2A_B_22_10(),
.F2A_B_22_11(),
.F2A_B_22_12(),
.F2A_B_22_13(),
.F2A_B_22_14(),
.F2A_B_22_15(),
.F2A_B_22_16(),
.F2A_B_22_17(),
.F2A_B_22_2(),
.F2A_B_22_3(),
.F2A_B_22_4(),
.F2A_B_22_5(),
.F2A_B_22_6(),
.F2A_B_22_7(),
.F2A_B_22_8(),
.F2A_B_22_9(),
.F2A_B_23_0(),
.F2A_B_23_1(),
.F2A_B_23_10(),
.F2A_B_23_11(),
.F2A_B_23_2(),
.F2A_B_23_3(),
.F2A_B_23_4(),
.F2A_B_23_5(),
.F2A_B_23_6(),
.F2A_B_23_7(),
.F2A_B_23_8(),
.F2A_B_23_9(),
.F2A_B_24_0(),
.F2A_B_24_1(),
.F2A_B_24_10(),
.F2A_B_24_11(),
.F2A_B_24_12(),
.F2A_B_24_13(),
.F2A_B_24_14(),
.F2A_B_24_15(),
.F2A_B_24_16(),
.F2A_B_24_17(),
.F2A_B_24_2(),
.F2A_B_24_3(),
.F2A_B_24_4(),
.F2A_B_24_5(),
.F2A_B_24_6(),
.F2A_B_24_7(),
.F2A_B_24_8(),
.F2A_B_24_9(),
.F2A_B_25_0(),
.F2A_B_25_1(),
.F2A_B_25_10(),
.F2A_B_25_11(),
.F2A_B_25_2(),
.F2A_B_25_3(),
.F2A_B_25_4(),
.F2A_B_25_5(),
.F2A_B_25_6(),
.F2A_B_25_7(),
.F2A_B_25_8(),
.F2A_B_25_9(),
.F2A_B_26_0(),
.F2A_B_26_1(),
.F2A_B_26_10(),
.F2A_B_26_11(),
.F2A_B_26_12(),
.F2A_B_26_13(),
.F2A_B_26_14(),
.F2A_B_26_15(),
.F2A_B_26_16(),
.F2A_B_26_17(),
.F2A_B_26_2(),
.F2A_B_26_3(),
.F2A_B_26_4(),
.F2A_B_26_5(),
.F2A_B_26_6(),
.F2A_B_26_7(),
.F2A_B_26_8(),
.F2A_B_26_9(),
.F2A_B_27_0(),
.F2A_B_27_1(),
.F2A_B_27_10(),
.F2A_B_27_11(),
.F2A_B_27_2(),
.F2A_B_27_3(),
.F2A_B_27_4(),
.F2A_B_27_5(),
.F2A_B_27_6(),
.F2A_B_27_7(),
.F2A_B_27_8(),
.F2A_B_27_9(),
.F2A_B_28_0(),
.F2A_B_28_1(),
.F2A_B_28_10(),
.F2A_B_28_11(),
.F2A_B_28_12(),
.F2A_B_28_13(),
.F2A_B_28_14(),
.F2A_B_28_15(),
.F2A_B_28_16(),
.F2A_B_28_17(),
.F2A_B_28_2(),
.F2A_B_28_3(),
.F2A_B_28_4(),
.F2A_B_28_5(),
.F2A_B_28_6(),
.F2A_B_28_7(),
.F2A_B_28_8(),
.F2A_B_28_9(),
.F2A_B_29_0(),
.F2A_B_29_1(),
.F2A_B_29_10(),
.F2A_B_29_11(),
.F2A_B_29_2(),
.F2A_B_29_3(),
.F2A_B_29_4(),
.F2A_B_29_5(),
.F2A_B_29_6(),
.F2A_B_29_7(),
.F2A_B_29_8(),
.F2A_B_29_9(),
.F2A_B_2_0(),
.F2A_B_2_1(),
.F2A_B_2_10(),
.F2A_B_2_11(),
.F2A_B_2_12(),
.F2A_B_2_13(),
.F2A_B_2_14(),
.F2A_B_2_15(),
.F2A_B_2_16(),
.F2A_B_2_17(),
.F2A_B_2_2(),
.F2A_B_2_3(),
.F2A_B_2_4(),
.F2A_B_2_5(),
.F2A_B_2_6(),
.F2A_B_2_7(),
.F2A_B_2_8(),
.F2A_B_2_9(),
.F2A_B_30_0(),
.F2A_B_30_1(),
.F2A_B_30_10(),
.F2A_B_30_11(),
.F2A_B_30_12(),
.F2A_B_30_13(),
.F2A_B_30_14(),
.F2A_B_30_15(),
.F2A_B_30_16(),
.F2A_B_30_17(),
.F2A_B_30_2(),
.F2A_B_30_3(),
.F2A_B_30_4(),
.F2A_B_30_5(),
.F2A_B_30_6(),
.F2A_B_30_7(),
.F2A_B_30_8(),
.F2A_B_30_9(),
.F2A_B_31_0(),
.F2A_B_31_1(),
.F2A_B_31_10(),
.F2A_B_31_11(),
.F2A_B_31_2(),
.F2A_B_31_3(),
.F2A_B_31_4(),
.F2A_B_31_5(),
.F2A_B_31_6(),
.F2A_B_31_7(),
.F2A_B_31_8(),
.F2A_B_31_9(),
.F2A_B_32_0(),
.F2A_B_32_1(),
.F2A_B_32_10(),
.F2A_B_32_11(),
.F2A_B_32_12(),
.F2A_B_32_13(),
.F2A_B_32_14(),
.F2A_B_32_15(),
.F2A_B_32_16(),
.F2A_B_32_17(),
.F2A_B_32_2(),
.F2A_B_32_3(),
.F2A_B_32_4(),
.F2A_B_32_5(),
.F2A_B_32_6(),
.F2A_B_32_7(),
.F2A_B_32_8(),
.F2A_B_32_9(),
.F2A_B_3_0(),
.F2A_B_3_1(),
.F2A_B_3_10(),
.F2A_B_3_11(),
.F2A_B_3_2(),
.F2A_B_3_3(),
.F2A_B_3_4(),
.F2A_B_3_5(),
.F2A_B_3_6(),
.F2A_B_3_7(),
.F2A_B_3_8(),
.F2A_B_3_9(),
.F2A_B_4_0(),
.F2A_B_4_1(),
.F2A_B_4_10(),
.F2A_B_4_11(),
.F2A_B_4_12(),
.F2A_B_4_13(),
.F2A_B_4_14(),
.F2A_B_4_15(),
.F2A_B_4_16(),
.F2A_B_4_17(),
.F2A_B_4_2(),
.F2A_B_4_3(),
.F2A_B_4_4(),
.F2A_B_4_5(),
.F2A_B_4_6(),
.F2A_B_4_7(),
.F2A_B_4_8(),
.F2A_B_4_9(),
.F2A_B_5_0(),
.F2A_B_5_1(),
.F2A_B_5_10(),
.F2A_B_5_11(),
.F2A_B_5_2(),
.F2A_B_5_3(),
.F2A_B_5_4(),
.F2A_B_5_5(),
.F2A_B_5_6(),
.F2A_B_5_7(),
.F2A_B_5_8(),
.F2A_B_5_9(),
.F2A_B_6_0(),
.F2A_B_6_1(),
.F2A_B_6_10(),
.F2A_B_6_11(),
.F2A_B_6_12(),
.F2A_B_6_13(),
.F2A_B_6_14(),
.F2A_B_6_15(),
.F2A_B_6_16(),
.F2A_B_6_17(),
.F2A_B_6_2(),
.F2A_B_6_3(),
.F2A_B_6_4(),
.F2A_B_6_5(),
.F2A_B_6_6(),
.F2A_B_6_7(),
.F2A_B_6_8(),
.F2A_B_6_9(),
.F2A_B_7_0(),
.F2A_B_7_1(),
.F2A_B_7_10(),
.F2A_B_7_11(),
.F2A_B_7_2(),
.F2A_B_7_3(),
.F2A_B_7_4(),
.F2A_B_7_5(),
.F2A_B_7_6(),
.F2A_B_7_7(),
.F2A_B_7_8(),
.F2A_B_7_9(),
.F2A_B_8_0(),
.F2A_B_8_1(),
.F2A_B_8_10(),
.F2A_B_8_11(),
.F2A_B_8_12(),
.F2A_B_8_13(),
.F2A_B_8_14(),
.F2A_B_8_15(),
.F2A_B_8_16(),
.F2A_B_8_17(),
.F2A_B_8_2(),
.F2A_B_8_3(),
.F2A_B_8_4(),
.F2A_B_8_5(),
.F2A_B_8_6(),
.F2A_B_8_7(),
.F2A_B_8_8(),
.F2A_B_8_9(),
.F2A_B_9_0(),
.F2A_B_9_1(),
.F2A_B_9_10(),
.F2A_B_9_11(),
.F2A_B_9_2(),
.F2A_B_9_3(),
.F2A_B_9_4(),
.F2A_B_9_5(),
.F2A_B_9_6(),
.F2A_B_9_7(),
.F2A_B_9_8(),
.F2A_B_9_9(),
.F2A_L_10_0(fpgaio_oe_20_o),
.F2A_L_10_1(fpgaio_data_20_o),
.F2A_L_10_10(fpgaio_oe_25_o),
.F2A_L_10_11(fpgaio_data_25_o),
.F2A_L_10_12(fpgaio_oe_26_o),
.F2A_L_10_13(fpgaio_data_26_o),
.F2A_L_10_14(fpgaio_oe_27_o),
.F2A_L_10_15(fpgaio_data_27_o),
.F2A_L_10_16(),
.F2A_L_10_17(),
.F2A_L_10_2(fpgaio_oe_21_o),
.F2A_L_10_3(fpgaio_data_21_o),
.F2A_L_10_4(fpgaio_oe_22_o),
.F2A_L_10_5(fpgaio_data_22_o),
.F2A_L_10_6(fpgaio_oe_23_o),
.F2A_L_10_7(fpgaio_data_23_o),
.F2A_L_10_8(fpgaio_oe_24_o),
.F2A_L_10_9(fpgaio_data_24_o),
.F2A_L_11_0(events_12_o),
.F2A_L_11_1(events_13_o),
.F2A_L_11_10(fpgaio_oe_19_o),
.F2A_L_11_11(fpgaio_data_19_o),
.F2A_L_11_2(events_14_o),
.F2A_L_11_3(events_15_o),
.F2A_L_11_4(fpgaio_oe_16_o),
.F2A_L_11_5(fpgaio_data_16_o),
.F2A_L_11_6(fpgaio_oe_17_o),
.F2A_L_11_7(fpgaio_data_17_o),
.F2A_L_11_8(fpgaio_oe_18_o),
.F2A_L_11_9(fpgaio_data_18_o),
.F2A_L_12_0(udma_cfg_data_26_o),
.F2A_L_12_1(udma_cfg_data_27_o),
.F2A_L_12_10(events_4_o),
.F2A_L_12_11(events_5_o),
.F2A_L_12_12(events_6_o),
.F2A_L_12_13(events_7_o),
.F2A_L_12_14(events_8_o),
.F2A_L_12_15(events_9_o),
.F2A_L_12_16(events_10_o),
.F2A_L_12_17(events_11_o),
.F2A_L_12_2(udma_cfg_data_28_o),
.F2A_L_12_3(udma_cfg_data_29_o),
.F2A_L_12_4(udma_cfg_data_30_o),
.F2A_L_12_5(udma_cfg_data_31_o),
.F2A_L_12_6(events_0_o),
.F2A_L_12_7(events_1_o),
.F2A_L_12_8(events_2_o),
.F2A_L_12_9(events_3_o),
.F2A_L_13_0(udma_cfg_data_14_o),
.F2A_L_13_1(udma_cfg_data_15_o),
.F2A_L_13_10(udma_cfg_data_24_o),
.F2A_L_13_11(udma_cfg_data_25_o),
.F2A_L_13_2(udma_cfg_data_16_o),
.F2A_L_13_3(udma_cfg_data_17_o),
.F2A_L_13_4(udma_cfg_data_18_o),
.F2A_L_13_5(udma_cfg_data_19_o),
.F2A_L_13_6(udma_cfg_data_20_o),
.F2A_L_13_7(udma_cfg_data_21_o),
.F2A_L_13_8(udma_cfg_data_22_o),
.F2A_L_13_9(udma_cfg_data_23_o),
.F2A_L_14_0(udma_rx_lin_data_28_o),
.F2A_L_14_1(udma_rx_lin_data_29_o),
.F2A_L_14_10(udma_cfg_data_6_o),
.F2A_L_14_11(udma_cfg_data_7_o),
.F2A_L_14_12(udma_cfg_data_8_o),
.F2A_L_14_13(udma_cfg_data_9_o),
.F2A_L_14_14(udma_cfg_data_10_o),
.F2A_L_14_15(udma_cfg_data_11_o),
.F2A_L_14_16(udma_cfg_data_12_o),
.F2A_L_14_17(udma_cfg_data_13_o),
.F2A_L_14_2(udma_rx_lin_data_30_o),
.F2A_L_14_3(udma_rx_lin_data_31_o),
.F2A_L_14_4(udma_cfg_data_0_o),
.F2A_L_14_5(udma_cfg_data_1_o),
.F2A_L_14_6(udma_cfg_data_2_o),
.F2A_L_14_7(udma_cfg_data_3_o),
.F2A_L_14_8(udma_cfg_data_4_o),
.F2A_L_14_9(udma_cfg_data_5_o),
.F2A_L_15_0(udma_rx_lin_data_16_o),
.F2A_L_15_1(udma_rx_lin_data_17_o),
.F2A_L_15_10(udma_rx_lin_data_26_o),
.F2A_L_15_11(udma_rx_lin_data_27_o),
.F2A_L_15_2(udma_rx_lin_data_18_o),
.F2A_L_15_3(udma_rx_lin_data_19_o),
.F2A_L_15_4(udma_rx_lin_data_20_o),
.F2A_L_15_5(udma_rx_lin_data_21_o),
.F2A_L_15_6(udma_rx_lin_data_22_o),
.F2A_L_15_7(udma_rx_lin_data_23_o),
.F2A_L_15_8(udma_rx_lin_data_24_o),
.F2A_L_15_9(udma_rx_lin_data_25_o),
.F2A_L_16_0(udma_tx_lin_ready_o),
.F2A_L_16_1(udma_rx_lin_valid_o),
.F2A_L_16_10(udma_rx_lin_data_8_o),
.F2A_L_16_11(udma_rx_lin_data_9_o),
.F2A_L_16_12(udma_rx_lin_data_10_o),
.F2A_L_16_13(udma_rx_lin_data_11_o),
.F2A_L_16_14(udma_rx_lin_data_12_o),
.F2A_L_16_15(udma_rx_lin_data_13_o),
.F2A_L_16_16(udma_rx_lin_data_14_o),
.F2A_L_16_17(udma_rx_lin_data_15_o),
.F2A_L_16_2(udma_rx_lin_data_0_o),
.F2A_L_16_3(udma_rx_lin_data_1_o),
.F2A_L_16_4(udma_rx_lin_data_2_o),
.F2A_L_16_5(udma_rx_lin_data_3_o),
.F2A_L_16_6(udma_rx_lin_data_4_o),
.F2A_L_16_7(udma_rx_lin_data_5_o),
.F2A_L_16_8(udma_rx_lin_data_6_o),
.F2A_L_16_9(udma_rx_lin_data_7_o),
.F2A_L_17_0(apb_hwce_prdata_0_o),
.F2A_L_17_1(apb_hwce_prdata_1_o),
.F2A_L_17_10(apb_hwce_prdata_10_o),
.F2A_L_17_11(apb_hwce_prdata_11_o),
.F2A_L_17_2(apb_hwce_prdata_2_o),
.F2A_L_17_3(apb_hwce_prdata_3_o),
.F2A_L_17_4(apb_hwce_prdata_4_o),
.F2A_L_17_5(apb_hwce_prdata_5_o),
.F2A_L_17_6(apb_hwce_prdata_6_o),
.F2A_L_17_7(apb_hwce_prdata_7_o),
.F2A_L_17_8(apb_hwce_prdata_8_o),
.F2A_L_17_9(apb_hwce_prdata_9_o),
.F2A_L_18_0(apb_hwce_prdata_12_o),
.F2A_L_18_1(apb_hwce_prdata_13_o),
.F2A_L_18_10(apb_hwce_prdata_22_o),
.F2A_L_18_11(apb_hwce_prdata_23_o),
.F2A_L_18_12(apb_hwce_prdata_24_o),
.F2A_L_18_13(apb_hwce_prdata_25_o),
.F2A_L_18_14(apb_hwce_prdata_26_o),
.F2A_L_18_15(apb_hwce_prdata_27_o),
.F2A_L_18_16(apb_hwce_prdata_28_o),
.F2A_L_18_17(apb_hwce_prdata_29_o),
.F2A_L_18_2(apb_hwce_prdata_14_o),
.F2A_L_18_3(apb_hwce_prdata_15_o),
.F2A_L_18_4(apb_hwce_prdata_16_o),
.F2A_L_18_5(apb_hwce_prdata_17_o),
.F2A_L_18_6(apb_hwce_prdata_18_o),
.F2A_L_18_7(apb_hwce_prdata_19_o),
.F2A_L_18_8(apb_hwce_prdata_20_o),
.F2A_L_18_9(apb_hwce_prdata_21_o),
.F2A_L_19_0(apb_hwce_prdata_30_o),
.F2A_L_19_1(apb_hwce_prdata_31_o),
.F2A_L_19_10(fpgaio_oe_31_o),
.F2A_L_19_11(fpgaio_data_31_o),
.F2A_L_19_2(apb_hwce_ready_o),
.F2A_L_19_3(apb_hwce_pslverr_o),
.F2A_L_19_4(fpgaio_oe_28_o),
.F2A_L_19_5(fpgaio_data_28_o),
.F2A_L_19_6(fpgaio_oe_29_o),
.F2A_L_19_7(fpgaio_data_29_o),
.F2A_L_19_8(fpgaio_oe_30_o),
.F2A_L_19_9(fpgaio_data_30_o),
.F2A_L_1_0(),
.F2A_L_1_1(),
.F2A_L_1_10(),
.F2A_L_1_11(),
.F2A_L_1_2(),
.F2A_L_1_3(),
.F2A_L_1_4(),
.F2A_L_1_5(),
.F2A_L_1_6(),
.F2A_L_1_7(),
.F2A_L_1_8(),
.F2A_L_1_9(),
.F2A_L_20_0(fpgaio_oe_32_o),
.F2A_L_20_1(fpgaio_data_32_o),
.F2A_L_20_10(fpgaio_oe_37_o),
.F2A_L_20_11(fpgaio_data_37_o),
.F2A_L_20_12(fpgaio_oe_38_o),
.F2A_L_20_13(fpgaio_data_38_o),
.F2A_L_20_14(fpgaio_oe_39_o),
.F2A_L_20_15(fpgaio_data_39_o),
.F2A_L_20_16(fpgaio_oe_40_o),
.F2A_L_20_17(fpgaio_data_40_o),
.F2A_L_20_2(fpgaio_oe_33_o),
.F2A_L_20_3(fpgaio_data_33_o),
.F2A_L_20_4(fpgaio_oe_34_o),
.F2A_L_20_5(fpgaio_data_34_o),
.F2A_L_20_6(fpgaio_oe_35_o),
.F2A_L_20_7(fpgaio_data_35_o),
.F2A_L_20_8(fpgaio_oe_36_o),
.F2A_L_20_9(fpgaio_data_36_o),
.F2A_L_21_0(fpgaio_oe_41_o),
.F2A_L_21_1(fpgaio_data_41_o),
.F2A_L_21_10(),
.F2A_L_21_11(),
.F2A_L_21_2(fpgaio_oe_42_o),
.F2A_L_21_3(fpgaio_data_42_o),
.F2A_L_21_4(),
.F2A_L_21_5(),
.F2A_L_21_6(),
.F2A_L_21_7(),
.F2A_L_21_8(),
.F2A_L_21_9(),
.F2A_L_22_0(),
.F2A_L_22_1(),
.F2A_L_22_10(),
.F2A_L_22_11(),
.F2A_L_22_12(),
.F2A_L_22_13(),
.F2A_L_22_14(),
.F2A_L_22_15(),
.F2A_L_22_16(),
.F2A_L_22_17(),
.F2A_L_22_2(),
.F2A_L_22_3(),
.F2A_L_22_4(),
.F2A_L_22_5(),
.F2A_L_22_6(),
.F2A_L_22_7(),
.F2A_L_22_8(),
.F2A_L_22_9(),
.F2A_L_23_0(),
.F2A_L_23_1(),
.F2A_L_23_10(),
.F2A_L_23_11(),
.F2A_L_23_2(),
.F2A_L_23_3(),
.F2A_L_23_4(),
.F2A_L_23_5(),
.F2A_L_23_6(),
.F2A_L_23_7(),
.F2A_L_23_8(),
.F2A_L_23_9(),
.F2A_L_24_0(),
.F2A_L_24_1(),
.F2A_L_24_10(),
.F2A_L_24_11(),
.F2A_L_24_12(),
.F2A_L_24_13(),
.F2A_L_24_14(),
.F2A_L_24_15(),
.F2A_L_24_16(),
.F2A_L_24_17(),
.F2A_L_24_2(),
.F2A_L_24_3(),
.F2A_L_24_4(),
.F2A_L_24_5(),
.F2A_L_24_6(),
.F2A_L_24_7(),
.F2A_L_24_8(),
.F2A_L_24_9(),
.F2A_L_25_0(),
.F2A_L_25_1(),
.F2A_L_25_10(),
.F2A_L_25_11(),
.F2A_L_25_2(),
.F2A_L_25_3(),
.F2A_L_25_4(),
.F2A_L_25_5(),
.F2A_L_25_6(),
.F2A_L_25_7(),
.F2A_L_25_8(),
.F2A_L_25_9(),
.F2A_L_26_0(),
.F2A_L_26_1(),
.F2A_L_26_10(),
.F2A_L_26_11(),
.F2A_L_26_12(),
.F2A_L_26_13(),
.F2A_L_26_14(),
.F2A_L_26_15(),
.F2A_L_26_16(),
.F2A_L_26_17(),
.F2A_L_26_2(),
.F2A_L_26_3(),
.F2A_L_26_4(),
.F2A_L_26_5(),
.F2A_L_26_6(),
.F2A_L_26_7(),
.F2A_L_26_8(),
.F2A_L_26_9(),
.F2A_L_27_0(),
.F2A_L_27_1(),
.F2A_L_27_10(),
.F2A_L_27_11(),
.F2A_L_27_2(),
.F2A_L_27_3(),
.F2A_L_27_4(),
.F2A_L_27_5(),
.F2A_L_27_6(),
.F2A_L_27_7(),
.F2A_L_27_8(),
.F2A_L_27_9(),
.F2A_L_28_0(),
.F2A_L_28_1(),
.F2A_L_28_10(),
.F2A_L_28_11(),
.F2A_L_28_12(),
.F2A_L_28_13(),
.F2A_L_28_14(),
.F2A_L_28_15(),
.F2A_L_28_16(),
.F2A_L_28_17(),
.F2A_L_28_2(),
.F2A_L_28_3(),
.F2A_L_28_4(),
.F2A_L_28_5(),
.F2A_L_28_6(),
.F2A_L_28_7(),
.F2A_L_28_8(),
.F2A_L_28_9(),
.F2A_L_29_0(),
.F2A_L_29_1(),
.F2A_L_29_10(),
.F2A_L_29_11(),
.F2A_L_29_2(),
.F2A_L_29_3(),
.F2A_L_29_4(),
.F2A_L_29_5(),
.F2A_L_29_6(),
.F2A_L_29_7(),
.F2A_L_29_8(),
.F2A_L_29_9(),
.F2A_L_2_0(),
.F2A_L_2_1(),
.F2A_L_2_10(),
.F2A_L_2_11(),
.F2A_L_2_12(),
.F2A_L_2_13(),
.F2A_L_2_14(),
.F2A_L_2_15(),
.F2A_L_2_16(),
.F2A_L_2_17(),
.F2A_L_2_2(),
.F2A_L_2_3(),
.F2A_L_2_4(),
.F2A_L_2_5(),
.F2A_L_2_6(),
.F2A_L_2_7(),
.F2A_L_2_8(),
.F2A_L_2_9(),
.F2A_L_30_0(),
.F2A_L_30_1(),
.F2A_L_30_10(),
.F2A_L_30_11(),
.F2A_L_30_12(),
.F2A_L_30_13(),
.F2A_L_30_14(),
.F2A_L_30_15(),
.F2A_L_30_16(),
.F2A_L_30_17(),
.F2A_L_30_2(),
.F2A_L_30_3(),
.F2A_L_30_4(),
.F2A_L_30_5(),
.F2A_L_30_6(),
.F2A_L_30_7(),
.F2A_L_30_8(),
.F2A_L_30_9(),
.F2A_L_31_0(),
.F2A_L_31_1(),
.F2A_L_31_10(),
.F2A_L_31_11(),
.F2A_L_31_2(),
.F2A_L_31_3(),
.F2A_L_31_4(),
.F2A_L_31_5(),
.F2A_L_31_6(),
.F2A_L_31_7(),
.F2A_L_31_8(),
.F2A_L_31_9(),
.F2A_L_32_0(),
.F2A_L_32_1(),
.F2A_L_32_10(),
.F2A_L_32_11(),
.F2A_L_32_12(),
.F2A_L_32_13(),
.F2A_L_32_14(),
.F2A_L_32_15(),
.F2A_L_32_16(),
.F2A_L_32_17(),
.F2A_L_32_2(),
.F2A_L_32_3(),
.F2A_L_32_4(),
.F2A_L_32_5(),
.F2A_L_32_6(),
.F2A_L_32_7(),
.F2A_L_32_8(),
.F2A_L_32_9(),
.F2A_L_3_0(),
.F2A_L_3_1(),
.F2A_L_3_10(),
.F2A_L_3_11(),
.F2A_L_3_2(),
.F2A_L_3_3(),
.F2A_L_3_4(),
.F2A_L_3_5(),
.F2A_L_3_6(),
.F2A_L_3_7(),
.F2A_L_3_8(),
.F2A_L_3_9(),
.F2A_L_4_0(),
.F2A_L_4_1(),
.F2A_L_4_10(),
.F2A_L_4_11(),
.F2A_L_4_12(),
.F2A_L_4_13(),
.F2A_L_4_14(),
.F2A_L_4_15(),
.F2A_L_4_16(),
.F2A_L_4_17(),
.F2A_L_4_2(),
.F2A_L_4_3(),
.F2A_L_4_4(),
.F2A_L_4_5(),
.F2A_L_4_6(),
.F2A_L_4_7(),
.F2A_L_4_8(),
.F2A_L_4_9(),
.F2A_L_5_0(),
.F2A_L_5_1(),
.F2A_L_5_10(),
.F2A_L_5_11(),
.F2A_L_5_2(),
.F2A_L_5_3(),
.F2A_L_5_4(),
.F2A_L_5_5(),
.F2A_L_5_6(),
.F2A_L_5_7(),
.F2A_L_5_8(),
.F2A_L_5_9(),
.F2A_L_6_0(),
.F2A_L_6_1(),
.F2A_L_6_10(),
.F2A_L_6_11(),
.F2A_L_6_12(),
.F2A_L_6_13(),
.F2A_L_6_14(),
.F2A_L_6_15(),
.F2A_L_6_16(),
.F2A_L_6_17(),
.F2A_L_6_2(),
.F2A_L_6_3(),
.F2A_L_6_4(),
.F2A_L_6_5(),
.F2A_L_6_6(),
.F2A_L_6_7(),
.F2A_L_6_8(),
.F2A_L_6_9(),
.F2A_L_7_0(),
.F2A_L_7_1(),
.F2A_L_7_10(),
.F2A_L_7_11(),
.F2A_L_7_2(),
.F2A_L_7_3(),
.F2A_L_7_4(),
.F2A_L_7_5(),
.F2A_L_7_6(),
.F2A_L_7_7(),
.F2A_L_7_8(),
.F2A_L_7_9(),
.F2A_L_8_0(),
.F2A_L_8_1(),
.F2A_L_8_10(),
.F2A_L_8_11(),
.F2A_L_8_12(),
.F2A_L_8_13(),
.F2A_L_8_14(),
.F2A_L_8_15(),
.F2A_L_8_16(),
.F2A_L_8_17(),
.F2A_L_8_2(),
.F2A_L_8_3(),
.F2A_L_8_4(),
.F2A_L_8_5(),
.F2A_L_8_6(),
.F2A_L_8_7(),
.F2A_L_8_8(),
.F2A_L_8_9(),
.F2A_L_9_0(),
.F2A_L_9_1(),
.F2A_L_9_10(),
.F2A_L_9_11(),
.F2A_L_9_2(),
.F2A_L_9_3(),
.F2A_L_9_4(),
.F2A_L_9_5(),
.F2A_L_9_6(),
.F2A_L_9_7(),
.F2A_L_9_8(),
.F2A_L_9_9(),
.F2A_R_10_0(tcdm_addr_p3_16_o),
.F2A_R_10_1(tcdm_wdata_p3_16_o),
.F2A_R_10_10(tcdm_wdata_p3_22_o),
.F2A_R_10_11(tcdm_wdata_p3_23_o),
.F2A_R_10_12(tcdm_wdata_p3_24_o),
.F2A_R_10_13(tcdm_wdata_p3_25_o),
.F2A_R_10_14(tcdm_wdata_p3_26_o),
.F2A_R_10_15(tcdm_wdata_p3_27_o),
.F2A_R_10_16(tcdm_wdata_p3_28_o),
.F2A_R_10_17(tcdm_wdata_p3_29_o),
.F2A_R_10_2(tcdm_addr_p3_17_o),
.F2A_R_10_3(tcdm_wdata_p3_17_o),
.F2A_R_10_4(tcdm_addr_p3_18_o),
.F2A_R_10_5(tcdm_wdata_p3_18_o),
.F2A_R_10_6(tcdm_addr_p3_19_o),
.F2A_R_10_7(tcdm_wdata_p3_19_o),
.F2A_R_10_8(tcdm_wdata_p3_20_o),
.F2A_R_10_9(tcdm_wdata_p3_21_o),
.F2A_R_11_0(tcdm_addr_p3_10_o),
.F2A_R_11_1(tcdm_wdata_p3_10_o),
.F2A_R_11_10(tcdm_addr_p3_15_o),
.F2A_R_11_11(tcdm_wdata_p3_15_o),
.F2A_R_11_2(tcdm_addr_p3_11_o),
.F2A_R_11_3(tcdm_wdata_p3_11_o),
.F2A_R_11_4(tcdm_addr_p3_12_o),
.F2A_R_11_5(tcdm_wdata_p3_12_o),
.F2A_R_11_6(tcdm_addr_p3_13_o),
.F2A_R_11_7(tcdm_wdata_p3_13_o),
.F2A_R_11_8(tcdm_addr_p3_14_o),
.F2A_R_11_9(tcdm_wdata_p3_14_o),
.F2A_R_12_0(tcdm_addr_p3_1_o),
.F2A_R_12_1(tcdm_wdata_p3_1_o),
.F2A_R_12_10(tcdm_addr_p3_6_o),
.F2A_R_12_11(tcdm_wdata_p3_6_o),
.F2A_R_12_12(tcdm_addr_p3_7_o),
.F2A_R_12_13(tcdm_wdata_p3_7_o),
.F2A_R_12_14(tcdm_addr_p3_8_o),
.F2A_R_12_15(tcdm_wdata_p3_8_o),
.F2A_R_12_16(tcdm_addr_p3_9_o),
.F2A_R_12_17(tcdm_wdata_p3_9_o),
.F2A_R_12_2(tcdm_addr_p3_2_o),
.F2A_R_12_3(tcdm_wdata_p3_2_o),
.F2A_R_12_4(tcdm_addr_p3_3_o),
.F2A_R_12_5(tcdm_wdata_p3_3_o),
.F2A_R_12_6(tcdm_addr_p3_4_o),
.F2A_R_12_7(tcdm_wdata_p3_4_o),
.F2A_R_12_8(tcdm_addr_p3_5_o),
.F2A_R_12_9(tcdm_wdata_p3_5_o),
.F2A_R_13_0(tcdm_wdata_p2_28_o),
.F2A_R_13_1(tcdm_wdata_p2_29_o),
.F2A_R_13_10(tcdm_addr_p3_0_o),
.F2A_R_13_11(tcdm_wdata_p3_0_o),
.F2A_R_13_2(tcdm_wdata_p2_30_o),
.F2A_R_13_3(tcdm_wdata_p2_31_o),
.F2A_R_13_4(tcdm_req_p2_o),
.F2A_R_13_5(tcdm_wen_p2_o),
.F2A_R_13_6(tcdm_be_p2_0_o),
.F2A_R_13_7(tcdm_be_p2_1_o),
.F2A_R_13_8(tcdm_be_p2_2_o),
.F2A_R_13_9(tcdm_be_p2_3_o),
.F2A_R_14_0(tcdm_addr_p2_15_o),
.F2A_R_14_1(tcdm_wdata_p2_15_o),
.F2A_R_14_10(tcdm_wdata_p2_20_o),
.F2A_R_14_11(tcdm_wdata_p2_21_o),
.F2A_R_14_12(tcdm_wdata_p2_22_o),
.F2A_R_14_13(tcdm_wdata_p2_23_o),
.F2A_R_14_14(tcdm_wdata_p2_24_o),
.F2A_R_14_15(tcdm_wdata_p2_25_o),
.F2A_R_14_16(tcdm_wdata_p2_26_o),
.F2A_R_14_17(tcdm_wdata_p2_27_o),
.F2A_R_14_2(tcdm_addr_p2_16_o),
.F2A_R_14_3(tcdm_wdata_p2_16_o),
.F2A_R_14_4(tcdm_addr_p2_17_o),
.F2A_R_14_5(tcdm_wdata_p2_17_o),
.F2A_R_14_6(tcdm_addr_p2_18_o),
.F2A_R_14_7(tcdm_wdata_p2_18_o),
.F2A_R_14_8(tcdm_addr_p2_19_o),
.F2A_R_14_9(tcdm_wdata_p2_19_o),
.F2A_R_15_0(tcdm_addr_p2_9_o),
.F2A_R_15_1(tcdm_wdata_p2_9_o),
.F2A_R_15_10(tcdm_addr_p2_14_o),
.F2A_R_15_11(tcdm_wdata_p2_14_o),
.F2A_R_15_2(tcdm_addr_p2_10_o),
.F2A_R_15_3(tcdm_wdata_p2_10_o),
.F2A_R_15_4(tcdm_addr_p2_11_o),
.F2A_R_15_5(tcdm_wdata_p2_11_o),
.F2A_R_15_6(tcdm_addr_p2_12_o),
.F2A_R_15_7(tcdm_wdata_p2_12_o),
.F2A_R_15_8(tcdm_addr_p2_13_o),
.F2A_R_15_9(tcdm_wdata_p2_13_o),
.F2A_R_16_0(tcdm_addr_p2_0_o),
.F2A_R_16_1(tcdm_wdata_p2_0_o),
.F2A_R_16_10(tcdm_addr_p2_5_o),
.F2A_R_16_11(tcdm_wdata_p2_5_o),
.F2A_R_16_12(tcdm_addr_p2_6_o),
.F2A_R_16_13(tcdm_wdata_p2_6_o),
.F2A_R_16_14(tcdm_addr_p2_7_o),
.F2A_R_16_15(tcdm_wdata_p2_7_o),
.F2A_R_16_16(tcdm_addr_p2_8_o),
.F2A_R_16_17(tcdm_wdata_p2_8_o),
.F2A_R_16_2(tcdm_addr_p2_1_o),
.F2A_R_16_3(tcdm_wdata_p2_1_o),
.F2A_R_16_4(tcdm_addr_p2_2_o),
.F2A_R_16_5(tcdm_wdata_p2_2_o),
.F2A_R_16_6(tcdm_addr_p2_3_o),
.F2A_R_16_7(tcdm_wdata_p2_3_o),
.F2A_R_16_8(tcdm_addr_p2_4_o),
.F2A_R_16_9(tcdm_wdata_p2_4_o),
.F2A_R_17_0(tcdm_addr_p0_0_o),
.F2A_R_17_1(tcdm_wdata_p0_0_o),
.F2A_R_17_10(tcdm_addr_p0_5_o),
.F2A_R_17_11(tcdm_wdata_p0_5_o),
.F2A_R_17_2(tcdm_addr_p0_1_o),
.F2A_R_17_3(tcdm_wdata_p0_1_o),
.F2A_R_17_4(tcdm_addr_p0_2_o),
.F2A_R_17_5(tcdm_wdata_p0_2_o),
.F2A_R_17_6(tcdm_addr_p0_3_o),
.F2A_R_17_7(tcdm_wdata_p0_3_o),
.F2A_R_17_8(tcdm_addr_p0_4_o),
.F2A_R_17_9(tcdm_wdata_p0_4_o),
.F2A_R_18_0(tcdm_addr_p0_6_o),
.F2A_R_18_1(tcdm_wdata_p0_6_o),
.F2A_R_18_10(tcdm_addr_p0_11_o),
.F2A_R_18_11(tcdm_wdata_p0_11_o),
.F2A_R_18_12(tcdm_addr_p0_12_o),
.F2A_R_18_13(tcdm_wdata_p0_12_o),
.F2A_R_18_14(tcdm_addr_p0_13_o),
.F2A_R_18_15(tcdm_wdata_p0_13_o),
.F2A_R_18_16(tcdm_addr_p0_14_o),
.F2A_R_18_17(tcdm_wdata_p0_14_o),
.F2A_R_18_2(tcdm_addr_p0_7_o),
.F2A_R_18_3(tcdm_wdata_p0_7_o),
.F2A_R_18_4(tcdm_addr_p0_8_o),
.F2A_R_18_5(tcdm_wdata_p0_8_o),
.F2A_R_18_6(tcdm_addr_p0_9_o),
.F2A_R_18_7(tcdm_wdata_p0_9_o),
.F2A_R_18_8(tcdm_addr_p0_10_o),
.F2A_R_18_9(tcdm_wdata_p0_10_o),
.F2A_R_19_0(tcdm_addr_p0_15_o),
.F2A_R_19_1(tcdm_wdata_p0_15_o),
.F2A_R_19_10(tcdm_wdata_p0_20_o),
.F2A_R_19_11(tcdm_wdata_p0_21_o),
.F2A_R_19_2(tcdm_addr_p0_16_o),
.F2A_R_19_3(tcdm_wdata_p0_16_o),
.F2A_R_19_4(tcdm_addr_p0_17_o),
.F2A_R_19_5(tcdm_wdata_p0_17_o),
.F2A_R_19_6(tcdm_addr_p0_18_o),
.F2A_R_19_7(tcdm_wdata_p0_18_o),
.F2A_R_19_8(tcdm_addr_p0_19_o),
.F2A_R_19_9(tcdm_wdata_p0_19_o),
.F2A_R_1_0(),
.F2A_R_1_1(),
.F2A_R_1_10(),
.F2A_R_1_11(),
.F2A_R_1_2(),
.F2A_R_1_3(),
.F2A_R_1_4(),
.F2A_R_1_5(),
.F2A_R_1_6(),
.F2A_R_1_7(),
.F2A_R_1_8(),
.F2A_R_1_9(),
.F2A_R_20_0(tcdm_wdata_p0_22_o),
.F2A_R_20_1(tcdm_wdata_p0_23_o),
.F2A_R_20_10(tcdm_req_p0_o),
.F2A_R_20_11(tcdm_wen_p0_o),
.F2A_R_20_12(tcdm_be_p0_0_o),
.F2A_R_20_13(tcdm_be_p0_1_o),
.F2A_R_20_14(tcdm_be_p0_2_o),
.F2A_R_20_15(tcdm_be_p0_3_o),
.F2A_R_20_16(tcdm_addr_p1_0_o),
.F2A_R_20_17(tcdm_wdata_p1_0_o),
.F2A_R_20_2(tcdm_wdata_p0_24_o),
.F2A_R_20_3(tcdm_wdata_p0_25_o),
.F2A_R_20_4(tcdm_wdata_p0_26_o),
.F2A_R_20_5(tcdm_wdata_p0_27_o),
.F2A_R_20_6(tcdm_wdata_p0_28_o),
.F2A_R_20_7(tcdm_wdata_p0_29_o),
.F2A_R_20_8(tcdm_wdata_p0_30_o),
.F2A_R_20_9(tcdm_wdata_p0_31_o),
.F2A_R_21_0(tcdm_addr_p1_1_o),
.F2A_R_21_1(tcdm_wdata_p1_1_o),
.F2A_R_21_10(tcdm_addr_p1_6_o),
.F2A_R_21_11(tcdm_wdata_p1_6_o),
.F2A_R_21_2(tcdm_addr_p1_2_o),
.F2A_R_21_3(tcdm_wdata_p1_2_o),
.F2A_R_21_4(tcdm_addr_p1_3_o),
.F2A_R_21_5(tcdm_wdata_p1_3_o),
.F2A_R_21_6(tcdm_addr_p1_4_o),
.F2A_R_21_7(tcdm_wdata_p1_4_o),
.F2A_R_21_8(tcdm_addr_p1_5_o),
.F2A_R_21_9(tcdm_wdata_p1_5_o),
.F2A_R_22_0(tcdm_addr_p1_7_o),
.F2A_R_22_1(tcdm_wdata_p1_7_o),
.F2A_R_22_10(tcdm_addr_p1_12_o),
.F2A_R_22_11(tcdm_wdata_p1_12_o),
.F2A_R_22_12(tcdm_addr_p1_13_o),
.F2A_R_22_13(tcdm_wdata_p1_13_o),
.F2A_R_22_14(tcdm_addr_p1_14_o),
.F2A_R_22_15(tcdm_wdata_p1_14_o),
.F2A_R_22_16(tcdm_addr_p1_15_o),
.F2A_R_22_17(tcdm_wdata_p1_15_o),
.F2A_R_22_2(tcdm_addr_p1_8_o),
.F2A_R_22_3(tcdm_wdata_p1_8_o),
.F2A_R_22_4(tcdm_addr_p1_9_o),
.F2A_R_22_5(tcdm_wdata_p1_9_o),
.F2A_R_22_6(tcdm_addr_p1_10_o),
.F2A_R_22_7(tcdm_wdata_p1_10_o),
.F2A_R_22_8(tcdm_addr_p1_11_o),
.F2A_R_22_9(tcdm_wdata_p1_11_o),
.F2A_R_23_0(tcdm_addr_p1_16_o),
.F2A_R_23_1(tcdm_wdata_p1_16_o),
.F2A_R_23_10(tcdm_wdata_p1_22_o),
.F2A_R_23_11(tcdm_wdata_p1_23_o),
.F2A_R_23_2(tcdm_addr_p1_17_o),
.F2A_R_23_3(tcdm_wdata_p1_17_o),
.F2A_R_23_4(tcdm_addr_p1_18_o),
.F2A_R_23_5(tcdm_wdata_p1_18_o),
.F2A_R_23_6(tcdm_addr_p1_19_o),
.F2A_R_23_7(tcdm_wdata_p1_19_o),
.F2A_R_23_8(tcdm_wdata_p1_20_o),
.F2A_R_23_9(tcdm_wdata_p1_21_o),
.F2A_R_24_0(tcdm_wdata_p1_24_o),
.F2A_R_24_1(tcdm_wdata_p1_25_o),
.F2A_R_24_10(tcdm_be_p1_0_o),
.F2A_R_24_11(tcdm_be_p1_1_o),
.F2A_R_24_12(tcdm_be_p1_2_o),
.F2A_R_24_13(tcdm_be_p1_3_o),
.F2A_R_24_14(fpgaio_oe_8_o),
.F2A_R_24_15(fpgaio_data_8_o),
.F2A_R_24_16(fpgaio_oe_9_o),
.F2A_R_24_17(fpgaio_data_9_o),
.F2A_R_24_2(tcdm_wdata_p1_26_o),
.F2A_R_24_3(tcdm_wdata_p1_27_o),
.F2A_R_24_4(tcdm_wdata_p1_28_o),
.F2A_R_24_5(tcdm_wdata_p1_29_o),
.F2A_R_24_6(tcdm_wdata_p1_30_o),
.F2A_R_24_7(tcdm_wdata_p1_31_o),
.F2A_R_24_8(tcdm_req_p1_o),
.F2A_R_24_9(tcdm_wen_p1_o),
.F2A_R_25_0(fpgaio_oe_10_o),
.F2A_R_25_1(fpgaio_data_10_o),
.F2A_R_25_10(),
.F2A_R_25_11(),
.F2A_R_25_2(fpgaio_oe_11_o),
.F2A_R_25_3(fpgaio_data_11_o),
.F2A_R_25_4(),
.F2A_R_25_5(),
.F2A_R_25_6(),
.F2A_R_25_7(),
.F2A_R_25_8(),
.F2A_R_25_9(),
.F2A_R_26_0(),
.F2A_R_26_1(),
.F2A_R_26_10(),
.F2A_R_26_11(),
.F2A_R_26_12(),
.F2A_R_26_13(),
.F2A_R_26_14(),
.F2A_R_26_15(),
.F2A_R_26_16(),
.F2A_R_26_17(),
.F2A_R_26_2(),
.F2A_R_26_3(),
.F2A_R_26_4(),
.F2A_R_26_5(),
.F2A_R_26_6(),
.F2A_R_26_7(),
.F2A_R_26_8(),
.F2A_R_26_9(),
.F2A_R_27_0(),
.F2A_R_27_1(),
.F2A_R_27_10(),
.F2A_R_27_11(),
.F2A_R_27_2(),
.F2A_R_27_3(),
.F2A_R_27_4(),
.F2A_R_27_5(),
.F2A_R_27_6(),
.F2A_R_27_7(),
.F2A_R_27_8(),
.F2A_R_27_9(),
.F2A_R_28_0(),
.F2A_R_28_1(),
.F2A_R_28_10(),
.F2A_R_28_11(),
.F2A_R_28_12(),
.F2A_R_28_13(),
.F2A_R_28_14(),
.F2A_R_28_15(),
.F2A_R_28_16(),
.F2A_R_28_17(),
.F2A_R_28_2(),
.F2A_R_28_3(),
.F2A_R_28_4(),
.F2A_R_28_5(),
.F2A_R_28_6(),
.F2A_R_28_7(),
.F2A_R_28_8(),
.F2A_R_28_9(),
.F2A_R_29_0(),
.F2A_R_29_1(),
.F2A_R_29_10(),
.F2A_R_29_11(),
.F2A_R_29_2(),
.F2A_R_29_3(),
.F2A_R_29_4(),
.F2A_R_29_5(),
.F2A_R_29_6(),
.F2A_R_29_7(),
.F2A_R_29_8(),
.F2A_R_29_9(),
.F2A_R_2_0(),
.F2A_R_2_1(),
.F2A_R_2_10(),
.F2A_R_2_11(),
.F2A_R_2_12(),
.F2A_R_2_13(),
.F2A_R_2_14(),
.F2A_R_2_15(),
.F2A_R_2_16(),
.F2A_R_2_17(),
.F2A_R_2_2(),
.F2A_R_2_3(),
.F2A_R_2_4(),
.F2A_R_2_5(),
.F2A_R_2_6(),
.F2A_R_2_7(),
.F2A_R_2_8(),
.F2A_R_2_9(),
.F2A_R_30_0(),
.F2A_R_30_1(),
.F2A_R_30_10(),
.F2A_R_30_11(),
.F2A_R_30_12(),
.F2A_R_30_13(),
.F2A_R_30_14(),
.F2A_R_30_15(),
.F2A_R_30_16(),
.F2A_R_30_17(),
.F2A_R_30_2(),
.F2A_R_30_3(),
.F2A_R_30_4(),
.F2A_R_30_5(),
.F2A_R_30_6(),
.F2A_R_30_7(),
.F2A_R_30_8(),
.F2A_R_30_9(),
.F2A_R_31_0(),
.F2A_R_31_1(),
.F2A_R_31_10(),
.F2A_R_31_11(),
.F2A_R_31_2(),
.F2A_R_31_3(),
.F2A_R_31_4(),
.F2A_R_31_5(),
.F2A_R_31_6(),
.F2A_R_31_7(),
.F2A_R_31_8(),
.F2A_R_31_9(),
.F2A_R_32_0(),
.F2A_R_32_1(),
.F2A_R_32_10(),
.F2A_R_32_11(),
.F2A_R_32_12(),
.F2A_R_32_13(),
.F2A_R_32_14(),
.F2A_R_32_15(),
.F2A_R_32_16(),
.F2A_R_32_17(),
.F2A_R_32_2(),
.F2A_R_32_3(),
.F2A_R_32_4(),
.F2A_R_32_5(),
.F2A_R_32_6(),
.F2A_R_32_7(),
.F2A_R_32_8(),
.F2A_R_32_9(),
.F2A_R_3_0(),
.F2A_R_3_1(),
.F2A_R_3_10(),
.F2A_R_3_11(),
.F2A_R_3_2(),
.F2A_R_3_3(),
.F2A_R_3_4(),
.F2A_R_3_5(),
.F2A_R_3_6(),
.F2A_R_3_7(),
.F2A_R_3_8(),
.F2A_R_3_9(),
.F2A_R_4_0(),
.F2A_R_4_1(),
.F2A_R_4_10(),
.F2A_R_4_11(),
.F2A_R_4_12(),
.F2A_R_4_13(),
.F2A_R_4_14(),
.F2A_R_4_15(),
.F2A_R_4_16(),
.F2A_R_4_17(),
.F2A_R_4_2(),
.F2A_R_4_3(),
.F2A_R_4_4(),
.F2A_R_4_5(),
.F2A_R_4_6(),
.F2A_R_4_7(),
.F2A_R_4_8(),
.F2A_R_4_9(),
.F2A_R_5_0(),
.F2A_R_5_1(),
.F2A_R_5_10(),
.F2A_R_5_11(),
.F2A_R_5_2(),
.F2A_R_5_3(),
.F2A_R_5_4(),
.F2A_R_5_5(),
.F2A_R_5_6(),
.F2A_R_5_7(),
.F2A_R_5_8(),
.F2A_R_5_9(),
.F2A_R_6_0(),
.F2A_R_6_1(),
.F2A_R_6_10(),
.F2A_R_6_11(),
.F2A_R_6_12(),
.F2A_R_6_13(),
.F2A_R_6_14(),
.F2A_R_6_15(),
.F2A_R_6_16(),
.F2A_R_6_17(),
.F2A_R_6_2(),
.F2A_R_6_3(),
.F2A_R_6_4(),
.F2A_R_6_5(),
.F2A_R_6_6(),
.F2A_R_6_7(),
.F2A_R_6_8(),
.F2A_R_6_9(),
.F2A_R_7_0(),
.F2A_R_7_1(),
.F2A_R_7_10(),
.F2A_R_7_11(),
.F2A_R_7_2(),
.F2A_R_7_3(),
.F2A_R_7_4(),
.F2A_R_7_5(),
.F2A_R_7_6(),
.F2A_R_7_7(),
.F2A_R_7_8(),
.F2A_R_7_9(),
.F2A_R_8_0(fpgaio_oe_14_o),
.F2A_R_8_1(fpgaio_data_14_o),
.F2A_R_8_10(),
.F2A_R_8_11(),
.F2A_R_8_12(),
.F2A_R_8_13(),
.F2A_R_8_14(),
.F2A_R_8_15(),
.F2A_R_8_16(),
.F2A_R_8_17(),
.F2A_R_8_2(fpgaio_oe_15_o),
.F2A_R_8_3(fpgaio_data_15_o),
.F2A_R_8_4(),
.F2A_R_8_5(),
.F2A_R_8_6(),
.F2A_R_8_7(),
.F2A_R_8_8(),
.F2A_R_8_9(),
.F2A_R_9_0(tcdm_wdata_p3_30_o),
.F2A_R_9_1(tcdm_wdata_p3_31_o),
.F2A_R_9_10(fpgaio_oe_13_o),
.F2A_R_9_11(fpgaio_data_13_o),
.F2A_R_9_2(tcdm_req_p3_o),
.F2A_R_9_3(tcdm_wen_p3_o),
.F2A_R_9_4(tcdm_be_p3_0_o),
.F2A_R_9_5(tcdm_be_p3_1_o),
.F2A_R_9_6(tcdm_be_p3_2_o),
.F2A_R_9_7(tcdm_be_p3_3_o),
.F2A_R_9_8(fpgaio_oe_12_o),
.F2A_R_9_9(fpgaio_data_12_o),
.F2A_T_10_0(MU0_EFPGA_MATHB_COEF_DATA_23_),
.F2A_T_10_1(MU0_EFPGA_MATHB_COEF_DATA_22_),
.F2A_T_10_10(MU0_EFPGA_MATHB_COEF_DATA_13_),
.F2A_T_10_11(MU0_EFPGA_MATHB_COEF_DATA_12_),
.F2A_T_10_12(MU0_EFPGA_MATHB_COEF_DATA_11_),
.F2A_T_10_13(MU0_EFPGA_MATHB_COEF_DATA_10_),
.F2A_T_10_14(MU0_EFPGA_MATHB_COEF_DATA_9_),
.F2A_T_10_15(MU0_EFPGA_MATHB_COEF_DATA_8_),
.F2A_T_10_16(MU0_EFPGA_MATHB_COEF_DATA_7_),
.F2A_T_10_17(MU0_EFPGA_MATHB_COEF_DATA_6_),
.F2A_T_10_2(MU0_EFPGA_MATHB_COEF_DATA_21_),
.F2A_T_10_3(MU0_EFPGA_MATHB_COEF_DATA_20_),
.F2A_T_10_4(MU0_EFPGA_MATHB_COEF_DATA_19_),
.F2A_T_10_5(MU0_EFPGA_MATHB_COEF_DATA_18_),
.F2A_T_10_6(MU0_EFPGA_MATHB_COEF_DATA_17_),
.F2A_T_10_7(MU0_EFPGA_MATHB_COEF_DATA_16_),
.F2A_T_10_8(MU0_EFPGA_MATHB_COEF_DATA_15_),
.F2A_T_10_9(MU0_EFPGA_MATHB_COEF_DATA_14_),
.F2A_T_11_0(MU0_EFPGA_MATHB_COEF_DATA_5_),
.F2A_T_11_1(MU0_EFPGA_MATHB_COEF_DATA_4_),
.F2A_T_11_10(MU0_EFPGA_TPRAM_COEF_W_DATA_31_),
.F2A_T_11_11(MU0_EFPGA_TPRAM_COEF_W_DATA_30_),
.F2A_T_11_2(MU0_EFPGA_MATHB_COEF_DATA_3_),
.F2A_T_11_3(MU0_EFPGA_MATHB_COEF_DATA_2_),
.F2A_T_11_4(MU0_EFPGA_MATHB_COEF_DATA_1_),
.F2A_T_11_5(MU0_EFPGA_MATHB_COEF_DATA_0_),
.F2A_T_11_6(MU0_EFPGA_MATHB_DATAOUT_SEL_1_),
.F2A_T_11_7(MU0_EFPGA_MATHB_DATAOUT_SEL_0_),
.F2A_T_11_8(MU0_EFPGA_TPRAM_COEF_W_MODE_1_),
.F2A_T_11_9(MU0_EFPGA_TPRAM_COEF_W_MODE_0_),
.F2A_T_12_0(MU0_EFPGA_TPRAM_COEF_W_DATA_29_),
.F2A_T_12_1(MU0_EFPGA_TPRAM_COEF_W_DATA_28_),
.F2A_T_12_10(MU0_EFPGA_TPRAM_COEF_W_DATA_19_),
.F2A_T_12_11(MU0_EFPGA_TPRAM_COEF_W_DATA_18_),
.F2A_T_12_12(MU0_EFPGA_TPRAM_COEF_W_DATA_17_),
.F2A_T_12_13(MU0_EFPGA_TPRAM_COEF_W_DATA_16_),
.F2A_T_12_14(MU0_EFPGA_TPRAM_COEF_W_DATA_15_),
.F2A_T_12_15(MU0_EFPGA_TPRAM_COEF_W_DATA_14_),
.F2A_T_12_16(MU0_EFPGA_TPRAM_COEF_W_DATA_13_),
.F2A_T_12_17(MU0_EFPGA_TPRAM_COEF_W_DATA_12_),
.F2A_T_12_2(MU0_EFPGA_TPRAM_COEF_W_DATA_27_),
.F2A_T_12_3(MU0_EFPGA_TPRAM_COEF_W_DATA_26_),
.F2A_T_12_4(MU0_EFPGA_TPRAM_COEF_W_DATA_25_),
.F2A_T_12_5(MU0_EFPGA_TPRAM_COEF_W_DATA_24_),
.F2A_T_12_6(MU0_EFPGA_TPRAM_COEF_W_DATA_23_),
.F2A_T_12_7(MU0_EFPGA_TPRAM_COEF_W_DATA_22_),
.F2A_T_12_8(MU0_EFPGA_TPRAM_COEF_W_DATA_21_),
.F2A_T_12_9(MU0_EFPGA_TPRAM_COEF_W_DATA_20_),
.F2A_T_13_0(MU0_EFPGA_TPRAM_COEF_W_DATA_11_),
.F2A_T_13_1(MU0_EFPGA_TPRAM_COEF_W_DATA_10_),
.F2A_T_13_10(MU0_EFPGA_TPRAM_COEF_W_DATA_1_),
.F2A_T_13_11(MU0_EFPGA_TPRAM_COEF_W_DATA_0_),
.F2A_T_13_2(MU0_EFPGA_TPRAM_COEF_W_DATA_9_),
.F2A_T_13_3(MU0_EFPGA_TPRAM_COEF_W_DATA_8_),
.F2A_T_13_4(MU0_EFPGA_TPRAM_COEF_W_DATA_7_),
.F2A_T_13_5(MU0_EFPGA_TPRAM_COEF_W_DATA_6_),
.F2A_T_13_6(MU0_EFPGA_TPRAM_COEF_W_DATA_5_),
.F2A_T_13_7(MU0_EFPGA_TPRAM_COEF_W_DATA_4_),
.F2A_T_13_8(MU0_EFPGA_TPRAM_COEF_W_DATA_3_),
.F2A_T_13_9(MU0_EFPGA_TPRAM_COEF_W_DATA_2_),
.F2A_T_14_0(MU0_EFPGA_TPRAM_COEF_W_CLK),
.F2A_T_14_1(MU0_EFPGA_TPRAM_COEF_W_ADDR_11_),
.F2A_T_14_10(MU0_EFPGA_TPRAM_COEF_W_ADDR_2_),
.F2A_T_14_11(MU0_EFPGA_TPRAM_COEF_W_ADDR_1_),
.F2A_T_14_12(MU0_EFPGA_TPRAM_COEF_W_ADDR_0_),
.F2A_T_14_13(MU0_EFPGA_TPRAM_COEF_WE),
.F2A_T_14_14(MU0_EFPGA_TPRAM_COEF_WDSEL),
.F2A_T_14_15(MU0_EFPGA_TPRAM_COEF_R_MODE_1_),
.F2A_T_14_16(MU0_EFPGA_TPRAM_COEF_R_MODE_0_),
.F2A_T_14_17(MU0_EFPGA_TPRAM_COEF_R_CLK),
.F2A_T_14_2(MU0_EFPGA_TPRAM_COEF_W_ADDR_10_),
.F2A_T_14_3(MU0_EFPGA_TPRAM_COEF_W_ADDR_9_),
.F2A_T_14_4(MU0_EFPGA_TPRAM_COEF_W_ADDR_8_),
.F2A_T_14_5(MU0_EFPGA_TPRAM_COEF_W_ADDR_7_),
.F2A_T_14_6(MU0_EFPGA_TPRAM_COEF_W_ADDR_6_),
.F2A_T_14_7(MU0_EFPGA_TPRAM_COEF_W_ADDR_5_),
.F2A_T_14_8(MU0_EFPGA_TPRAM_COEF_W_ADDR_4_),
.F2A_T_14_9(MU0_EFPGA_TPRAM_COEF_W_ADDR_3_),
.F2A_T_15_0(MU0_EFPGA_TPRAM_COEF_R_ADDR_11_),
.F2A_T_15_1(MU0_EFPGA_TPRAM_COEF_R_ADDR_10_),
.F2A_T_15_10(MU0_EFPGA_TPRAM_COEF_R_ADDR_1_),
.F2A_T_15_11(MU0_EFPGA_TPRAM_COEF_R_ADDR_0_),
.F2A_T_15_2(MU0_EFPGA_TPRAM_COEF_R_ADDR_9_),
.F2A_T_15_3(MU0_EFPGA_TPRAM_COEF_R_ADDR_8_),
.F2A_T_15_4(MU0_EFPGA_TPRAM_COEF_R_ADDR_7_),
.F2A_T_15_5(MU0_EFPGA_TPRAM_COEF_R_ADDR_6_),
.F2A_T_15_6(MU0_EFPGA_TPRAM_COEF_R_ADDR_5_),
.F2A_T_15_7(MU0_EFPGA_TPRAM_COEF_R_ADDR_4_),
.F2A_T_15_8(MU0_EFPGA_TPRAM_COEF_R_ADDR_3_),
.F2A_T_15_9(MU0_EFPGA_TPRAM_COEF_R_ADDR_2_),
.F2A_T_16_0(MU0_EFPGA_TPRAM_COEF_POWERDN),
.F2A_T_16_1(),
.F2A_T_16_10(),
.F2A_T_16_11(),
.F2A_T_16_12(),
.F2A_T_16_13(),
.F2A_T_16_17(),
.F2A_T_16_2(),
.F2A_T_16_3(),
.F2A_T_16_4(),
.F2A_T_16_5(),
.F2A_T_16_6(),
.F2A_T_16_7(),
.F2A_T_16_8(),
.F2A_T_16_9(),
.F2A_T_17_0(MU1_EFPGA_TPRAM_OPER_W_MODE_1_),
.F2A_T_17_1(MU1_EFPGA_TPRAM_OPER_W_MODE_0_),
.F2A_T_17_10(MU1_EFPGA_TPRAM_OPER_W_DATA_23_),
.F2A_T_17_11(MU1_EFPGA_TPRAM_OPER_W_DATA_22_),
.F2A_T_17_2(MU1_EFPGA_TPRAM_OPER_W_DATA_31_),
.F2A_T_17_3(MU1_EFPGA_TPRAM_OPER_W_DATA_30_),
.F2A_T_17_4(MU1_EFPGA_TPRAM_OPER_W_DATA_29_),
.F2A_T_17_5(MU1_EFPGA_TPRAM_OPER_W_DATA_28_),
.F2A_T_17_6(MU1_EFPGA_TPRAM_OPER_W_DATA_27_),
.F2A_T_17_7(MU1_EFPGA_TPRAM_OPER_W_DATA_26_),
.F2A_T_17_8(MU1_EFPGA_TPRAM_OPER_W_DATA_25_),
.F2A_T_17_9(MU1_EFPGA_TPRAM_OPER_W_DATA_24_),
.F2A_T_18_0(MU1_EFPGA_TPRAM_OPER_W_DATA_21_),
.F2A_T_18_1(MU1_EFPGA_TPRAM_OPER_W_DATA_20_),
.F2A_T_18_10(MU1_EFPGA_TPRAM_OPER_W_DATA_11_),
.F2A_T_18_11(MU1_EFPGA_TPRAM_OPER_W_DATA_10_),
.F2A_T_18_12(MU1_EFPGA_TPRAM_OPER_W_DATA_9_),
.F2A_T_18_13(MU1_EFPGA_TPRAM_OPER_W_DATA_8_),
.F2A_T_18_14(MU1_EFPGA_TPRAM_OPER_W_DATA_7_),
.F2A_T_18_15(MU1_EFPGA_TPRAM_OPER_W_DATA_6_),
.F2A_T_18_16(MU1_EFPGA_TPRAM_OPER_W_DATA_5_),
.F2A_T_18_17(MU1_EFPGA_TPRAM_OPER_W_DATA_4_),
.F2A_T_18_2(MU1_EFPGA_TPRAM_OPER_W_DATA_19_),
.F2A_T_18_3(MU1_EFPGA_TPRAM_OPER_W_DATA_18_),
.F2A_T_18_4(MU1_EFPGA_TPRAM_OPER_W_DATA_17_),
.F2A_T_18_5(MU1_EFPGA_TPRAM_OPER_W_DATA_16_),
.F2A_T_18_6(MU1_EFPGA_TPRAM_OPER_W_DATA_15_),
.F2A_T_18_7(MU1_EFPGA_TPRAM_OPER_W_DATA_14_),
.F2A_T_18_8(MU1_EFPGA_TPRAM_OPER_W_DATA_13_),
.F2A_T_18_9(MU1_EFPGA_TPRAM_OPER_W_DATA_12_),
.F2A_T_19_0(MU1_EFPGA_TPRAM_OPER_W_DATA_3_),
.F2A_T_19_1(MU1_EFPGA_TPRAM_OPER_W_DATA_2_),
.F2A_T_19_10(MU1_EFPGA_TPRAM_OPER_W_ADDR_6_),
.F2A_T_19_11(MU1_EFPGA_TPRAM_OPER_W_ADDR_5_),
.F2A_T_19_2(MU1_EFPGA_TPRAM_OPER_W_DATA_1_),
.F2A_T_19_3(MU1_EFPGA_TPRAM_OPER_W_DATA_0_),
.F2A_T_19_4(MU1_EFPGA_TPRAM_OPER_W_CLK),
.F2A_T_19_5(MU1_EFPGA_TPRAM_OPER_W_ADDR_11_),
.F2A_T_19_6(MU1_EFPGA_TPRAM_OPER_W_ADDR_10_),
.F2A_T_19_7(MU1_EFPGA_TPRAM_OPER_W_ADDR_9_),
.F2A_T_19_8(MU1_EFPGA_TPRAM_OPER_W_ADDR_8_),
.F2A_T_19_9(MU1_EFPGA_TPRAM_OPER_W_ADDR_7_),
.F2A_T_1_0(),
.F2A_T_1_1(),
.F2A_T_1_10(),
.F2A_T_1_11(),
.F2A_T_1_2(),
.F2A_T_1_3(),
.F2A_T_1_4(),
.F2A_T_1_5(),
.F2A_T_1_6(),
.F2A_T_1_7(),
.F2A_T_1_8(),
.F2A_T_1_9(),
.F2A_T_20_0(MU1_EFPGA_TPRAM_OPER_W_ADDR_4_),
.F2A_T_20_1(MU1_EFPGA_TPRAM_OPER_W_ADDR_3_),
.F2A_T_20_10(MU1_EFPGA_TPRAM_OPER_R_ADDR_11_),
.F2A_T_20_11(MU1_EFPGA_TPRAM_OPER_R_ADDR_10_),
.F2A_T_20_12(MU1_EFPGA_TPRAM_OPER_R_ADDR_9_),
.F2A_T_20_13(MU1_EFPGA_TPRAM_OPER_R_ADDR_8_),
.F2A_T_20_14(MU1_EFPGA_TPRAM_OPER_R_ADDR_7_),
.F2A_T_20_15(MU1_EFPGA_TPRAM_OPER_R_ADDR_6_),
.F2A_T_20_16(MU1_EFPGA_TPRAM_OPER_R_ADDR_5_),
.F2A_T_20_17(MU1_EFPGA_TPRAM_OPER_R_ADDR_4_),
.F2A_T_20_2(MU1_EFPGA_TPRAM_OPER_W_ADDR_2_),
.F2A_T_20_3(MU1_EFPGA_TPRAM_OPER_W_ADDR_1_),
.F2A_T_20_4(MU1_EFPGA_TPRAM_OPER_W_ADDR_0_),
.F2A_T_20_5(MU1_EFPGA_TPRAM_OPER_WE),
.F2A_T_20_6(MU1_EFPGA_TPRAM_OPER_WDSEL),
.F2A_T_20_7(MU1_EFPGA_TPRAM_OPER_R_MODE_1_),
.F2A_T_20_8(MU1_EFPGA_TPRAM_OPER_R_MODE_0_),
.F2A_T_20_9(MU1_EFPGA_TPRAM_OPER_R_CLK),
.F2A_T_21_0(MU1_EFPGA_TPRAM_OPER_R_ADDR_3_),
.F2A_T_21_1(MU1_EFPGA_TPRAM_OPER_R_ADDR_2_),
.F2A_T_21_10(MU1_EFPGA_MATHB_MAC_OUT_SEL_2_),
.F2A_T_21_11(MU1_EFPGA_MATHB_MAC_OUT_SEL_1_),
.F2A_T_21_2(MU1_EFPGA_TPRAM_OPER_R_ADDR_1_),
.F2A_T_21_3(MU1_EFPGA_TPRAM_OPER_R_ADDR_0_),
.F2A_T_21_4(MU1_EFPGA_TPRAM_OPER_POWERDN),
.F2A_T_21_5(MU1_EFPGA2MATHB_CLK),
.F2A_T_21_6(MU1_EFPGA_MATHB_CLK_EN),
.F2A_T_21_7(MU1_EFPGA_MATHB_MAC_OUT_SEL_5_),
.F2A_T_21_8(MU1_EFPGA_MATHB_MAC_OUT_SEL_4_),
.F2A_T_21_9(MU1_EFPGA_MATHB_MAC_OUT_SEL_3_),
.F2A_T_22_0(MU1_EFPGA_MATHB_MAC_OUT_SEL_0_),
.F2A_T_22_1(MU1_EFPGA_MATHB_MAC_ACC_SAT),
.F2A_T_22_10(MU1_EFPGA_MATHB_OPER_DATA_26_),
.F2A_T_22_11(MU1_EFPGA_MATHB_OPER_DATA_25_),
.F2A_T_22_12(MU1_EFPGA_MATHB_OPER_DATA_24_),
.F2A_T_22_13(MU1_EFPGA_MATHB_OPER_DATA_23_),
.F2A_T_22_14(MU1_EFPGA_MATHB_OPER_DATA_22_),
.F2A_T_22_15(MU1_EFPGA_MATHB_OPER_DATA_21_),
.F2A_T_22_16(MU1_EFPGA_MATHB_OPER_DATA_20_),
.F2A_T_22_17(MU1_EFPGA_MATHB_OPER_DATA_19_),
.F2A_T_22_2(MU1_EFPGA_MATHB_MAC_ACC_RND),
.F2A_T_22_3(MU1_EFPGA_MATHB_MAC_ACC_CLEAR),
.F2A_T_22_4(MU1_EFPGA_MATHB_OPER_SEL),
.F2A_T_22_5(MU1_EFPGA_MATHB_OPER_DATA_31_),
.F2A_T_22_6(MU1_EFPGA_MATHB_OPER_DATA_30_),
.F2A_T_22_7(MU1_EFPGA_MATHB_OPER_DATA_29_),
.F2A_T_22_8(MU1_EFPGA_MATHB_OPER_DATA_28_),
.F2A_T_22_9(MU1_EFPGA_MATHB_OPER_DATA_27_),
.F2A_T_23_0(MU1_EFPGA_MATHB_OPER_DATA_18_),
.F2A_T_23_1(MU1_EFPGA_MATHB_OPER_DATA_17_),
.F2A_T_23_10(MU1_EFPGA_MATHB_OPER_DATA_8_),
.F2A_T_23_11(MU1_EFPGA_MATHB_OPER_DATA_7_),
.F2A_T_23_2(MU1_EFPGA_MATHB_OPER_DATA_16_),
.F2A_T_23_3(MU1_EFPGA_MATHB_OPER_DATA_15_),
.F2A_T_23_4(MU1_EFPGA_MATHB_OPER_DATA_14_),
.F2A_T_23_5(MU1_EFPGA_MATHB_OPER_DATA_13_),
.F2A_T_23_6(MU1_EFPGA_MATHB_OPER_DATA_12_),
.F2A_T_23_7(MU1_EFPGA_MATHB_OPER_DATA_11_),
.F2A_T_23_8(MU1_EFPGA_MATHB_OPER_DATA_10_),
.F2A_T_23_9(MU1_EFPGA_MATHB_OPER_DATA_9_),
.F2A_T_24_0(MU1_EFPGA_MATHB_OPER_DATA_6_),
.F2A_T_24_1(MU1_EFPGA_MATHB_OPER_DATA_5_),
.F2A_T_24_10(MU1_EFPGA_MATHB_COEF_DATA_29_),
.F2A_T_24_11(MU1_EFPGA_MATHB_COEF_DATA_28_),
.F2A_T_24_12(MU1_EFPGA_MATHB_COEF_DATA_27_),
.F2A_T_24_13(MU1_EFPGA_MATHB_COEF_DATA_26_),
.F2A_T_24_14(MU1_EFPGA_MATHB_COEF_DATA_25_),
.F2A_T_24_15(MU1_EFPGA_MATHB_COEF_DATA_24_),
.F2A_T_24_16(MU1_EFPGA_MATHB_COEF_DATA_23_),
.F2A_T_24_17(MU1_EFPGA_MATHB_COEF_DATA_22_),
.F2A_T_24_2(MU1_EFPGA_MATHB_OPER_DATA_4_),
.F2A_T_24_3(MU1_EFPGA_MATHB_OPER_DATA_3_),
.F2A_T_24_4(MU1_EFPGA_MATHB_OPER_DATA_2_),
.F2A_T_24_5(MU1_EFPGA_MATHB_OPER_DATA_1_),
.F2A_T_24_6(MU1_EFPGA_MATHB_OPER_DATA_0_),
.F2A_T_24_7(MU1_EFPGA_MATHB_COEF_SEL),
.F2A_T_24_8(MU1_EFPGA_MATHB_COEF_DATA_31_),
.F2A_T_24_9(MU1_EFPGA_MATHB_COEF_DATA_30_),
.F2A_T_25_0(MU1_EFPGA_MATHB_COEF_DATA_21_),
.F2A_T_25_1(MU1_EFPGA_MATHB_COEF_DATA_20_),
.F2A_T_25_10(MU1_EFPGA_MATHB_COEF_DATA_11_),
.F2A_T_25_11(MU1_EFPGA_MATHB_COEF_DATA_10_),
.F2A_T_25_2(MU1_EFPGA_MATHB_COEF_DATA_19_),
.F2A_T_25_3(MU1_EFPGA_MATHB_COEF_DATA_18_),
.F2A_T_25_4(MU1_EFPGA_MATHB_COEF_DATA_17_),
.F2A_T_25_5(MU1_EFPGA_MATHB_COEF_DATA_16_),
.F2A_T_25_6(MU1_EFPGA_MATHB_COEF_DATA_15_),
.F2A_T_25_7(MU1_EFPGA_MATHB_COEF_DATA_14_),
.F2A_T_25_8(MU1_EFPGA_MATHB_COEF_DATA_13_),
.F2A_T_25_9(MU1_EFPGA_MATHB_COEF_DATA_12_),
.F2A_T_26_0(MU1_EFPGA_MATHB_COEF_DATA_9_),
.F2A_T_26_1(MU1_EFPGA_MATHB_COEF_DATA_8_),
.F2A_T_26_10(MU1_EFPGA_MATHB_DATAOUT_SEL_1_),
.F2A_T_26_11(MU1_EFPGA_MATHB_DATAOUT_SEL_0_),
.F2A_T_26_12(MU1_EFPGA_TPRAM_COEF_W_MODE_1_),
.F2A_T_26_13(MU1_EFPGA_TPRAM_COEF_W_MODE_0_),
.F2A_T_26_14(MU1_EFPGA_TPRAM_COEF_W_DATA_31_),
.F2A_T_26_15(MU1_EFPGA_TPRAM_COEF_W_DATA_30_),
.F2A_T_26_16(MU1_EFPGA_TPRAM_COEF_W_DATA_29_),
.F2A_T_26_17(MU1_EFPGA_TPRAM_COEF_W_DATA_28_),
.F2A_T_26_2(MU1_EFPGA_MATHB_COEF_DATA_7_),
.F2A_T_26_3(MU1_EFPGA_MATHB_COEF_DATA_6_),
.F2A_T_26_4(MU1_EFPGA_MATHB_COEF_DATA_5_),
.F2A_T_26_5(MU1_EFPGA_MATHB_COEF_DATA_4_),
.F2A_T_26_6(MU1_EFPGA_MATHB_COEF_DATA_3_),
.F2A_T_26_7(MU1_EFPGA_MATHB_COEF_DATA_2_),
.F2A_T_26_8(MU1_EFPGA_MATHB_COEF_DATA_1_),
.F2A_T_26_9(MU1_EFPGA_MATHB_COEF_DATA_0_),
.F2A_T_27_0(MU1_EFPGA_TPRAM_COEF_W_DATA_27_),
.F2A_T_27_1(MU1_EFPGA_TPRAM_COEF_W_DATA_26_),
.F2A_T_27_10(MU1_EFPGA_TPRAM_COEF_W_DATA_17_),
.F2A_T_27_11(MU1_EFPGA_TPRAM_COEF_W_DATA_16_),
.F2A_T_27_2(MU1_EFPGA_TPRAM_COEF_W_DATA_25_),
.F2A_T_27_3(MU1_EFPGA_TPRAM_COEF_W_DATA_24_),
.F2A_T_27_4(MU1_EFPGA_TPRAM_COEF_W_DATA_23_),
.F2A_T_27_5(MU1_EFPGA_TPRAM_COEF_W_DATA_22_),
.F2A_T_27_6(MU1_EFPGA_TPRAM_COEF_W_DATA_21_),
.F2A_T_27_7(MU1_EFPGA_TPRAM_COEF_W_DATA_20_),
.F2A_T_27_8(MU1_EFPGA_TPRAM_COEF_W_DATA_19_),
.F2A_T_27_9(MU1_EFPGA_TPRAM_COEF_W_DATA_18_),
.F2A_T_28_0(MU1_EFPGA_TPRAM_COEF_W_DATA_15_),
.F2A_T_28_1(MU1_EFPGA_TPRAM_COEF_W_DATA_14_),
.F2A_T_28_10(MU1_EFPGA_TPRAM_COEF_W_DATA_5_),
.F2A_T_28_11(MU1_EFPGA_TPRAM_COEF_W_DATA_4_),
.F2A_T_28_12(MU1_EFPGA_TPRAM_COEF_W_DATA_3_),
.F2A_T_28_13(MU1_EFPGA_TPRAM_COEF_W_DATA_2_),
.F2A_T_28_14(MU1_EFPGA_TPRAM_COEF_W_DATA_1_),
.F2A_T_28_15(MU1_EFPGA_TPRAM_COEF_W_DATA_0_),
.F2A_T_28_16(MU1_EFPGA_TPRAM_COEF_W_CLK),
.F2A_T_28_17(MU1_EFPGA_TPRAM_COEF_W_ADDR_11_),
.F2A_T_28_2(MU1_EFPGA_TPRAM_COEF_W_DATA_13_),
.F2A_T_28_3(MU1_EFPGA_TPRAM_COEF_W_DATA_12_),
.F2A_T_28_4(MU1_EFPGA_TPRAM_COEF_W_DATA_11_),
.F2A_T_28_5(MU1_EFPGA_TPRAM_COEF_W_DATA_10_),
.F2A_T_28_6(MU1_EFPGA_TPRAM_COEF_W_DATA_9_),
.F2A_T_28_7(MU1_EFPGA_TPRAM_COEF_W_DATA_8_),
.F2A_T_28_8(MU1_EFPGA_TPRAM_COEF_W_DATA_7_),
.F2A_T_28_9(MU1_EFPGA_TPRAM_COEF_W_DATA_6_),
.F2A_T_29_0(MU1_EFPGA_TPRAM_COEF_W_ADDR_10_),
.F2A_T_29_1(MU1_EFPGA_TPRAM_COEF_W_ADDR_9_),
.F2A_T_29_10(MU1_EFPGA_TPRAM_COEF_W_ADDR_0_),
.F2A_T_29_11(MU1_EFPGA_TPRAM_COEF_WE),
.F2A_T_29_2(MU1_EFPGA_TPRAM_COEF_W_ADDR_8_),
.F2A_T_29_3(MU1_EFPGA_TPRAM_COEF_W_ADDR_7_),
.F2A_T_29_4(MU1_EFPGA_TPRAM_COEF_W_ADDR_6_),
.F2A_T_29_5(MU1_EFPGA_TPRAM_COEF_W_ADDR_5_),
.F2A_T_29_6(MU1_EFPGA_TPRAM_COEF_W_ADDR_4_),
.F2A_T_29_7(MU1_EFPGA_TPRAM_COEF_W_ADDR_3_),
.F2A_T_29_8(MU1_EFPGA_TPRAM_COEF_W_ADDR_2_),
.F2A_T_29_9(MU1_EFPGA_TPRAM_COEF_W_ADDR_1_),
.F2A_T_2_0(),
.F2A_T_2_1(),
.F2A_T_2_10(MU0_EFPGA_TPRAM_OPER_W_DATA_25_),
.F2A_T_2_11(MU0_EFPGA_TPRAM_OPER_W_DATA_24_),
.F2A_T_2_12(MU0_EFPGA_TPRAM_OPER_W_DATA_23_),
.F2A_T_2_13(MU0_EFPGA_TPRAM_OPER_W_DATA_22_),
.F2A_T_2_14(MU0_EFPGA_TPRAM_OPER_W_DATA_21_),
.F2A_T_2_15(MU0_EFPGA_TPRAM_OPER_W_DATA_20_),
.F2A_T_2_16(MU0_EFPGA_TPRAM_OPER_W_DATA_19_),
.F2A_T_2_17(MU0_EFPGA_TPRAM_OPER_W_DATA_18_),
.F2A_T_2_2(MU0_EFPGA_TPRAM_OPER_W_MODE_1_),
.F2A_T_2_3(MU0_EFPGA_TPRAM_OPER_W_MODE_0_),
.F2A_T_2_4(MU0_EFPGA_TPRAM_OPER_W_DATA_31_),
.F2A_T_2_5(MU0_EFPGA_TPRAM_OPER_W_DATA_30_),
.F2A_T_2_6(MU0_EFPGA_TPRAM_OPER_W_DATA_29_),
.F2A_T_2_7(MU0_EFPGA_TPRAM_OPER_W_DATA_28_),
.F2A_T_2_8(MU0_EFPGA_TPRAM_OPER_W_DATA_27_),
.F2A_T_2_9(MU0_EFPGA_TPRAM_OPER_W_DATA_26_),
.F2A_T_30_0(MU1_EFPGA_TPRAM_COEF_WDSEL),
.F2A_T_30_1(MU1_EFPGA_TPRAM_COEF_R_MODE_1_),
.F2A_T_30_10(MU1_EFPGA_TPRAM_COEF_R_ADDR_5_),
.F2A_T_30_11(MU1_EFPGA_TPRAM_COEF_R_ADDR_4_),
.F2A_T_30_12(MU1_EFPGA_TPRAM_COEF_R_ADDR_3_),
.F2A_T_30_13(MU1_EFPGA_TPRAM_COEF_R_ADDR_2_),
.F2A_T_30_14(MU1_EFPGA_TPRAM_COEF_R_ADDR_1_),
.F2A_T_30_15(MU1_EFPGA_TPRAM_COEF_R_ADDR_0_),
.F2A_T_30_16(MU1_EFPGA_TPRAM_COEF_POWERDN),
.F2A_T_30_17(),
.F2A_T_30_2(MU1_EFPGA_TPRAM_COEF_R_MODE_0_),
.F2A_T_30_3(MU1_EFPGA_TPRAM_COEF_R_CLK),
.F2A_T_30_4(MU1_EFPGA_TPRAM_COEF_R_ADDR_11_),
.F2A_T_30_5(MU1_EFPGA_TPRAM_COEF_R_ADDR_10_),
.F2A_T_30_6(MU1_EFPGA_TPRAM_COEF_R_ADDR_9_),
.F2A_T_30_7(MU1_EFPGA_TPRAM_COEF_R_ADDR_8_),
.F2A_T_30_8(MU1_EFPGA_TPRAM_COEF_R_ADDR_7_),
.F2A_T_30_9(MU1_EFPGA_TPRAM_COEF_R_ADDR_6_),
.F2A_T_31_0(),
.F2A_T_31_1(),
.F2A_T_31_10(),
.F2A_T_31_11(),
.F2A_T_31_2(),
.F2A_T_31_3(),
.F2A_T_31_4(),
.F2A_T_31_5(),
.F2A_T_31_6(),
.F2A_T_31_7(),
.F2A_T_31_8(),
.F2A_T_31_9(),
.F2A_T_32_0(),
.F2A_T_32_1(),
.F2A_T_32_10(),
.F2A_T_32_11(),
.F2A_T_32_12(),
.F2A_T_32_13(),
.F2A_T_32_14(),
.F2A_T_32_15(),
.F2A_T_32_16(),
.F2A_T_32_17(),
.F2A_T_32_2(),
.F2A_T_32_3(),
.F2A_T_32_4(),
.F2A_T_32_5(),
.F2A_T_32_6(),
.F2A_T_32_7(),
.F2A_T_32_8(),
.F2A_T_32_9(),
.F2A_T_3_0(MU0_EFPGA_TPRAM_OPER_W_DATA_17_),
.F2A_T_3_1(MU0_EFPGA_TPRAM_OPER_W_DATA_16_),
.F2A_T_3_10(MU0_EFPGA_TPRAM_OPER_W_DATA_7_),
.F2A_T_3_11(MU0_EFPGA_TPRAM_OPER_W_DATA_6_),
.F2A_T_3_2(MU0_EFPGA_TPRAM_OPER_W_DATA_15_),
.F2A_T_3_3(MU0_EFPGA_TPRAM_OPER_W_DATA_14_),
.F2A_T_3_4(MU0_EFPGA_TPRAM_OPER_W_DATA_13_),
.F2A_T_3_5(MU0_EFPGA_TPRAM_OPER_W_DATA_12_),
.F2A_T_3_6(MU0_EFPGA_TPRAM_OPER_W_DATA_11_),
.F2A_T_3_7(MU0_EFPGA_TPRAM_OPER_W_DATA_10_),
.F2A_T_3_8(MU0_EFPGA_TPRAM_OPER_W_DATA_9_),
.F2A_T_3_9(MU0_EFPGA_TPRAM_OPER_W_DATA_8_),
.F2A_T_4_0(MU0_EFPGA_TPRAM_OPER_W_DATA_5_),
.F2A_T_4_1(MU0_EFPGA_TPRAM_OPER_W_DATA_4_),
.F2A_T_4_10(MU0_EFPGA_TPRAM_OPER_W_ADDR_8_),
.F2A_T_4_11(MU0_EFPGA_TPRAM_OPER_W_ADDR_7_),
.F2A_T_4_12(MU0_EFPGA_TPRAM_OPER_W_ADDR_6_),
.F2A_T_4_13(MU0_EFPGA_TPRAM_OPER_W_ADDR_5_),
.F2A_T_4_14(MU0_EFPGA_TPRAM_OPER_W_ADDR_4_),
.F2A_T_4_15(MU0_EFPGA_TPRAM_OPER_W_ADDR_3_),
.F2A_T_4_16(MU0_EFPGA_TPRAM_OPER_W_ADDR_2_),
.F2A_T_4_17(MU0_EFPGA_TPRAM_OPER_W_ADDR_1_),
.F2A_T_4_2(MU0_EFPGA_TPRAM_OPER_W_DATA_3_),
.F2A_T_4_3(MU0_EFPGA_TPRAM_OPER_W_DATA_2_),
.F2A_T_4_4(MU0_EFPGA_TPRAM_OPER_W_DATA_1_),
.F2A_T_4_5(MU0_EFPGA_TPRAM_OPER_W_DATA_0_),
.F2A_T_4_6(MU0_EFPGA_TPRAM_OPER_W_CLK),
.F2A_T_4_7(MU0_EFPGA_TPRAM_OPER_W_ADDR_11_),
.F2A_T_4_8(MU0_EFPGA_TPRAM_OPER_W_ADDR_10_),
.F2A_T_4_9(MU0_EFPGA_TPRAM_OPER_W_ADDR_9_),
.F2A_T_5_0(MU0_EFPGA_TPRAM_OPER_W_ADDR_0_),
.F2A_T_5_1(MU0_EFPGA_TPRAM_OPER_WE),
.F2A_T_5_10(MU0_EFPGA_TPRAM_OPER_R_ADDR_7_),
.F2A_T_5_11(MU0_EFPGA_TPRAM_OPER_R_ADDR_6_),
.F2A_T_5_2(MU0_EFPGA_TPRAM_OPER_WDSEL),
.F2A_T_5_3(MU0_EFPGA_TPRAM_OPER_R_MODE_1_),
.F2A_T_5_4(MU0_EFPGA_TPRAM_OPER_R_MODE_0_),
.F2A_T_5_5(MU0_EFPGA_TPRAM_OPER_R_CLK),
.F2A_T_5_6(MU0_EFPGA_TPRAM_OPER_R_ADDR_11_),
.F2A_T_5_7(MU0_EFPGA_TPRAM_OPER_R_ADDR_10_),
.F2A_T_5_8(MU0_EFPGA_TPRAM_OPER_R_ADDR_9_),
.F2A_T_5_9(MU0_EFPGA_TPRAM_OPER_R_ADDR_8_),
.F2A_T_6_0(MU0_EFPGA_TPRAM_OPER_R_ADDR_5_),
.F2A_T_6_1(MU0_EFPGA_TPRAM_OPER_R_ADDR_4_),
.F2A_T_6_10(MU0_EFPGA_MATHB_MAC_OUT_SEL_4_),
.F2A_T_6_11(MU0_EFPGA_MATHB_MAC_OUT_SEL_3_),
.F2A_T_6_12(MU0_EFPGA_MATHB_MAC_OUT_SEL_2_),
.F2A_T_6_13(MU0_EFPGA_MATHB_MAC_OUT_SEL_1_),
.F2A_T_6_14(MU0_EFPGA_MATHB_MAC_OUT_SEL_0_),
.F2A_T_6_15(MU0_EFPGA_MATHB_MAC_ACC_SAT),
.F2A_T_6_16(MU0_EFPGA_MATHB_MAC_ACC_RND),
.F2A_T_6_17(MU0_EFPGA_MATHB_MAC_ACC_CLEAR),
.F2A_T_6_2(MU0_EFPGA_TPRAM_OPER_R_ADDR_3_),
.F2A_T_6_3(MU0_EFPGA_TPRAM_OPER_R_ADDR_2_),
.F2A_T_6_4(MU0_EFPGA_TPRAM_OPER_R_ADDR_1_),
.F2A_T_6_5(MU0_EFPGA_TPRAM_OPER_R_ADDR_0_),
.F2A_T_6_6(MU0_EFPGA_TPRAM_OPER_POWERDN),
.F2A_T_6_7(MU0_EFPGA2MATHB_CLK),
.F2A_T_6_8(MU0_EFPGA_MATHB_CLK_EN),
.F2A_T_6_9(MU0_EFPGA_MATHB_MAC_OUT_SEL_5_),
.F2A_T_7_0(MU0_EFPGA_MATHB_OPER_SEL),
.F2A_T_7_1(MU0_EFPGA_MATHB_OPER_DATA_31_),
.F2A_T_7_10(MU0_EFPGA_MATHB_OPER_DATA_22_),
.F2A_T_7_11(MU0_EFPGA_MATHB_OPER_DATA_21_),
.F2A_T_7_2(MU0_EFPGA_MATHB_OPER_DATA_30_),
.F2A_T_7_3(MU0_EFPGA_MATHB_OPER_DATA_29_),
.F2A_T_7_4(MU0_EFPGA_MATHB_OPER_DATA_28_),
.F2A_T_7_5(MU0_EFPGA_MATHB_OPER_DATA_27_),
.F2A_T_7_6(MU0_EFPGA_MATHB_OPER_DATA_26_),
.F2A_T_7_7(MU0_EFPGA_MATHB_OPER_DATA_25_),
.F2A_T_7_8(MU0_EFPGA_MATHB_OPER_DATA_24_),
.F2A_T_7_9(MU0_EFPGA_MATHB_OPER_DATA_23_),
.F2A_T_8_0(MU0_EFPGA_MATHB_OPER_DATA_20_),
.F2A_T_8_1(MU0_EFPGA_MATHB_OPER_DATA_19_),
.F2A_T_8_10(MU0_EFPGA_MATHB_OPER_DATA_10_),
.F2A_T_8_11(MU0_EFPGA_MATHB_OPER_DATA_9_),
.F2A_T_8_12(MU0_EFPGA_MATHB_OPER_DATA_8_),
.F2A_T_8_13(MU0_EFPGA_MATHB_OPER_DATA_7_),
.F2A_T_8_14(MU0_EFPGA_MATHB_OPER_DATA_6_),
.F2A_T_8_15(MU0_EFPGA_MATHB_OPER_DATA_5_),
.F2A_T_8_16(MU0_EFPGA_MATHB_OPER_DATA_4_),
.F2A_T_8_17(MU0_EFPGA_MATHB_OPER_DATA_3_),
.F2A_T_8_2(MU0_EFPGA_MATHB_OPER_DATA_18_),
.F2A_T_8_3(MU0_EFPGA_MATHB_OPER_DATA_17_),
.F2A_T_8_4(MU0_EFPGA_MATHB_OPER_DATA_16_),
.F2A_T_8_5(MU0_EFPGA_MATHB_OPER_DATA_15_),
.F2A_T_8_6(MU0_EFPGA_MATHB_OPER_DATA_14_),
.F2A_T_8_7(MU0_EFPGA_MATHB_OPER_DATA_13_),
.F2A_T_8_8(MU0_EFPGA_MATHB_OPER_DATA_12_),
.F2A_T_8_9(MU0_EFPGA_MATHB_OPER_DATA_11_),
.F2A_T_9_0(MU0_EFPGA_MATHB_OPER_DATA_2_),
.F2A_T_9_1(MU0_EFPGA_MATHB_OPER_DATA_1_),
.F2A_T_9_10(MU0_EFPGA_MATHB_COEF_DATA_25_),
.F2A_T_9_11(MU0_EFPGA_MATHB_COEF_DATA_24_),
.F2A_T_9_2(MU0_EFPGA_MATHB_OPER_DATA_0_),
.F2A_T_9_3(MU0_EFPGA_MATHB_COEF_SEL),
.F2A_T_9_4(MU0_EFPGA_MATHB_COEF_DATA_31_),
.F2A_T_9_5(MU0_EFPGA_MATHB_COEF_DATA_30_),
.F2A_T_9_6(MU0_EFPGA_MATHB_COEF_DATA_29_),
.F2A_T_9_7(MU0_EFPGA_MATHB_COEF_DATA_28_),
.F2A_T_9_8(MU0_EFPGA_MATHB_COEF_DATA_27_),
.F2A_T_9_9(MU0_EFPGA_MATHB_COEF_DATA_26_),
.F2Adef_B_10_0(),
.F2Adef_B_10_1(),
.F2Adef_B_10_2(),
.F2Adef_B_10_3(),
.F2Adef_B_10_4(),
.F2Adef_B_10_5(),
.F2Adef_B_10_6(),
.F2Adef_B_11_0(),
.F2Adef_B_11_1(),
.F2Adef_B_11_2(),
.F2Adef_B_11_3(),
.F2Adef_B_12_0(),
.F2Adef_B_12_1(),
.F2Adef_B_12_2(),
.F2Adef_B_12_3(),
.F2Adef_B_12_4(),
.F2Adef_B_12_5(),
.F2Adef_B_12_6(),
.F2Adef_B_13_0(),
.F2Adef_B_13_1(),
.F2Adef_B_13_2(),
.F2Adef_B_13_3(),
.F2Adef_B_14_0(),
.F2Adef_B_14_1(),
.F2Adef_B_14_2(),
.F2Adef_B_14_3(),
.F2Adef_B_14_4(),
.F2Adef_B_14_5(),
.F2Adef_B_14_6(),
.F2Adef_B_15_0(),
.F2Adef_B_15_1(),
.F2Adef_B_15_2(),
.F2Adef_B_15_3(),
.F2Adef_B_16_0(),
.F2Adef_B_16_1(),
.F2Adef_B_16_2(),
.F2Adef_B_16_3(),
.F2Adef_B_16_4(),
.F2Adef_B_16_5(),
.F2Adef_B_16_6(),
.F2Adef_B_17_0(),
.F2Adef_B_17_1(),
.F2Adef_B_17_2(),
.F2Adef_B_17_3(),
.F2Adef_B_18_0(),
.F2Adef_B_18_1(),
.F2Adef_B_18_2(),
.F2Adef_B_18_3(),
.F2Adef_B_18_4(),
.F2Adef_B_18_5(),
.F2Adef_B_18_6(),
.F2Adef_B_19_0(),
.F2Adef_B_19_1(),
.F2Adef_B_19_2(),
.F2Adef_B_19_3(),
.F2Adef_B_1_0(),
.F2Adef_B_1_1(),
.F2Adef_B_1_2(),
.F2Adef_B_1_3(),
.F2Adef_B_20_0(),
.F2Adef_B_20_1(),
.F2Adef_B_20_2(),
.F2Adef_B_20_3(),
.F2Adef_B_20_4(),
.F2Adef_B_20_5(),
.F2Adef_B_20_6(),
.F2Adef_B_21_0(),
.F2Adef_B_21_1(),
.F2Adef_B_21_2(),
.F2Adef_B_21_3(),
.F2Adef_B_22_0(),
.F2Adef_B_22_1(),
.F2Adef_B_22_2(),
.F2Adef_B_22_3(),
.F2Adef_B_22_4(),
.F2Adef_B_22_5(),
.F2Adef_B_22_6(),
.F2Adef_B_23_0(),
.F2Adef_B_23_1(),
.F2Adef_B_23_2(),
.F2Adef_B_23_3(),
.F2Adef_B_24_0(),
.F2Adef_B_24_1(),
.F2Adef_B_24_2(),
.F2Adef_B_24_3(),
.F2Adef_B_24_4(),
.F2Adef_B_24_5(),
.F2Adef_B_24_6(),
.F2Adef_B_25_0(),
.F2Adef_B_25_1(),
.F2Adef_B_25_2(),
.F2Adef_B_25_3(),
.F2Adef_B_26_0(),
.F2Adef_B_26_1(),
.F2Adef_B_26_2(),
.F2Adef_B_26_3(),
.F2Adef_B_26_4(),
.F2Adef_B_26_5(),
.F2Adef_B_26_6(),
.F2Adef_B_27_0(),
.F2Adef_B_27_1(),
.F2Adef_B_27_2(),
.F2Adef_B_27_3(),
.F2Adef_B_28_0(),
.F2Adef_B_28_1(),
.F2Adef_B_28_2(),
.F2Adef_B_28_3(),
.F2Adef_B_28_4(),
.F2Adef_B_28_5(),
.F2Adef_B_28_6(),
.F2Adef_B_29_0(),
.F2Adef_B_29_1(),
.F2Adef_B_29_2(),
.F2Adef_B_29_3(),
.F2Adef_B_2_0(),
.F2Adef_B_2_1(),
.F2Adef_B_2_2(),
.F2Adef_B_2_3(),
.F2Adef_B_2_4(),
.F2Adef_B_2_5(),
.F2Adef_B_2_6(),
.F2Adef_B_30_0(),
.F2Adef_B_30_1(),
.F2Adef_B_30_2(),
.F2Adef_B_30_3(),
.F2Adef_B_30_4(),
.F2Adef_B_30_5(),
.F2Adef_B_30_6(),
.F2Adef_B_31_0(),
.F2Adef_B_31_1(),
.F2Adef_B_31_2(),
.F2Adef_B_31_3(),
.F2Adef_B_32_0(),
.F2Adef_B_32_1(),
.F2Adef_B_32_2(),
.F2Adef_B_32_3(),
.F2Adef_B_32_4(),
.F2Adef_B_32_5(),
.F2Adef_B_32_6(),
.F2Adef_B_3_0(),
.F2Adef_B_3_1(),
.F2Adef_B_3_2(),
.F2Adef_B_3_3(),
.F2Adef_B_4_0(),
.F2Adef_B_4_1(),
.F2Adef_B_4_2(),
.F2Adef_B_4_3(),
.F2Adef_B_4_4(),
.F2Adef_B_4_5(),
.F2Adef_B_4_6(),
.F2Adef_B_5_0(),
.F2Adef_B_5_1(),
.F2Adef_B_5_2(),
.F2Adef_B_5_3(),
.F2Adef_B_6_0(),
.F2Adef_B_6_1(),
.F2Adef_B_6_2(),
.F2Adef_B_6_3(),
.F2Adef_B_6_4(),
.F2Adef_B_6_5(),
.F2Adef_B_6_6(),
.F2Adef_B_7_0(),
.F2Adef_B_7_1(),
.F2Adef_B_7_2(),
.F2Adef_B_7_3(),
.F2Adef_B_8_0(),
.F2Adef_B_8_1(),
.F2Adef_B_8_2(),
.F2Adef_B_8_3(),
.F2Adef_B_8_4(),
.F2Adef_B_8_5(),
.F2Adef_B_8_6(),
.F2Adef_B_9_0(),
.F2Adef_B_9_1(),
.F2Adef_B_9_2(),
.F2Adef_B_9_3(),
.F2Adef_L_10_0(),
.F2Adef_L_10_1(),
.F2Adef_L_10_2(),
.F2Adef_L_10_3(),
.F2Adef_L_10_4(),
.F2Adef_L_10_5(),
.F2Adef_L_10_6(),
.F2Adef_L_11_0(),
.F2Adef_L_11_1(),
.F2Adef_L_11_2(),
.F2Adef_L_11_3(),
.F2Adef_L_12_0(),
.F2Adef_L_12_1(),
.F2Adef_L_12_2(),
.F2Adef_L_12_3(),
.F2Adef_L_12_4(),
.F2Adef_L_12_5(),
.F2Adef_L_12_6(),
.F2Adef_L_13_0(),
.F2Adef_L_13_1(),
.F2Adef_L_13_2(),
.F2Adef_L_13_3(),
.F2Adef_L_14_0(),
.F2Adef_L_14_1(),
.F2Adef_L_14_2(),
.F2Adef_L_14_3(),
.F2Adef_L_14_4(),
.F2Adef_L_14_5(),
.F2Adef_L_14_6(),
.F2Adef_L_15_0(),
.F2Adef_L_15_1(),
.F2Adef_L_15_2(),
.F2Adef_L_15_3(),
.F2Adef_L_16_0(),
.F2Adef_L_16_1(),
.F2Adef_L_16_2(),
.F2Adef_L_16_3(),
.F2Adef_L_16_4(),
.F2Adef_L_16_5(),
.F2Adef_L_16_6(),
.F2Adef_L_17_0(),
.F2Adef_L_17_1(),
.F2Adef_L_17_2(),
.F2Adef_L_17_3(),
.F2Adef_L_18_0(),
.F2Adef_L_18_1(),
.F2Adef_L_18_2(),
.F2Adef_L_18_3(),
.F2Adef_L_18_4(),
.F2Adef_L_18_5(),
.F2Adef_L_18_6(),
.F2Adef_L_19_0(),
.F2Adef_L_19_1(),
.F2Adef_L_19_2(),
.F2Adef_L_19_3(),
.F2Adef_L_1_0(),
.F2Adef_L_1_1(),
.F2Adef_L_1_2(),
.F2Adef_L_1_3(),
.F2Adef_L_20_0(),
.F2Adef_L_20_1(),
.F2Adef_L_20_2(),
.F2Adef_L_20_3(),
.F2Adef_L_20_4(),
.F2Adef_L_20_5(),
.F2Adef_L_20_6(),
.F2Adef_L_21_0(),
.F2Adef_L_21_1(),
.F2Adef_L_21_2(),
.F2Adef_L_21_3(),
.F2Adef_L_22_0(),
.F2Adef_L_22_1(),
.F2Adef_L_22_2(),
.F2Adef_L_22_3(),
.F2Adef_L_22_4(),
.F2Adef_L_22_5(),
.F2Adef_L_22_6(),
.F2Adef_L_23_0(),
.F2Adef_L_23_1(),
.F2Adef_L_23_2(),
.F2Adef_L_23_3(),
.F2Adef_L_24_0(),
.F2Adef_L_24_1(),
.F2Adef_L_24_2(),
.F2Adef_L_24_3(),
.F2Adef_L_24_4(),
.F2Adef_L_24_5(),
.F2Adef_L_24_6(),
.F2Adef_L_25_0(),
.F2Adef_L_25_1(),
.F2Adef_L_25_2(),
.F2Adef_L_25_3(),
.F2Adef_L_26_0(),
.F2Adef_L_26_1(),
.F2Adef_L_26_2(),
.F2Adef_L_26_3(),
.F2Adef_L_26_4(),
.F2Adef_L_26_5(),
.F2Adef_L_26_6(),
.F2Adef_L_27_0(),
.F2Adef_L_27_1(),
.F2Adef_L_27_2(),
.F2Adef_L_27_3(),
.F2Adef_L_28_0(),
.F2Adef_L_28_1(),
.F2Adef_L_28_2(),
.F2Adef_L_28_3(),
.F2Adef_L_28_4(),
.F2Adef_L_28_5(),
.F2Adef_L_28_6(),
.F2Adef_L_29_0(),
.F2Adef_L_29_1(),
.F2Adef_L_29_2(),
.F2Adef_L_29_3(),
.F2Adef_L_2_0(),
.F2Adef_L_2_1(),
.F2Adef_L_2_2(),
.F2Adef_L_2_3(),
.F2Adef_L_2_4(),
.F2Adef_L_2_5(),
.F2Adef_L_2_6(),
.F2Adef_L_30_0(),
.F2Adef_L_30_1(),
.F2Adef_L_30_2(),
.F2Adef_L_30_3(),
.F2Adef_L_30_4(),
.F2Adef_L_30_5(),
.F2Adef_L_30_6(),
.F2Adef_L_31_0(),
.F2Adef_L_31_1(),
.F2Adef_L_31_2(),
.F2Adef_L_31_3(),
.F2Adef_L_32_0(),
.F2Adef_L_32_1(),
.F2Adef_L_32_2(),
.F2Adef_L_32_3(),
.F2Adef_L_32_4(),
.F2Adef_L_32_5(),
.F2Adef_L_32_6(),
.F2Adef_L_3_0(),
.F2Adef_L_3_1(),
.F2Adef_L_3_2(),
.F2Adef_L_3_3(),
.F2Adef_L_4_0(),
.F2Adef_L_4_1(),
.F2Adef_L_4_2(),
.F2Adef_L_4_3(),
.F2Adef_L_4_4(),
.F2Adef_L_4_5(),
.F2Adef_L_4_6(),
.F2Adef_L_5_0(),
.F2Adef_L_5_1(),
.F2Adef_L_5_2(),
.F2Adef_L_5_3(),
.F2Adef_L_6_0(),
.F2Adef_L_6_1(),
.F2Adef_L_6_2(),
.F2Adef_L_6_3(),
.F2Adef_L_6_4(),
.F2Adef_L_6_5(),
.F2Adef_L_6_6(),
.F2Adef_L_7_0(),
.F2Adef_L_7_1(),
.F2Adef_L_7_2(),
.F2Adef_L_7_3(),
.F2Adef_L_8_0(),
.F2Adef_L_8_1(),
.F2Adef_L_8_2(),
.F2Adef_L_8_3(),
.F2Adef_L_8_4(),
.F2Adef_L_8_5(),
.F2Adef_L_8_6(),
.F2Adef_L_9_0(),
.F2Adef_L_9_1(),
.F2Adef_L_9_2(),
.F2Adef_L_9_3(),
.F2Adef_R_10_0(),
.F2Adef_R_10_1(),
.F2Adef_R_10_2(),
.F2Adef_R_10_3(),
.F2Adef_R_10_4(),
.F2Adef_R_10_5(),
.F2Adef_R_10_6(),
.F2Adef_R_11_0(),
.F2Adef_R_11_1(),
.F2Adef_R_11_2(),
.F2Adef_R_11_3(),
.F2Adef_R_12_0(),
.F2Adef_R_12_1(),
.F2Adef_R_12_2(),
.F2Adef_R_12_3(),
.F2Adef_R_12_4(),
.F2Adef_R_12_5(),
.F2Adef_R_12_6(),
.F2Adef_R_13_0(),
.F2Adef_R_13_1(),
.F2Adef_R_13_2(),
.F2Adef_R_13_3(),
.F2Adef_R_14_0(),
.F2Adef_R_14_1(),
.F2Adef_R_14_2(),
.F2Adef_R_14_3(),
.F2Adef_R_14_4(),
.F2Adef_R_14_5(),
.F2Adef_R_14_6(),
.F2Adef_R_15_0(),
.F2Adef_R_15_1(),
.F2Adef_R_15_2(),
.F2Adef_R_15_3(),
.F2Adef_R_16_0(),
.F2Adef_R_16_1(),
.F2Adef_R_16_2(),
.F2Adef_R_16_3(),
.F2Adef_R_16_4(),
.F2Adef_R_16_5(),
.F2Adef_R_16_6(),
.F2Adef_R_17_0(),
.F2Adef_R_17_1(),
.F2Adef_R_17_2(),
.F2Adef_R_17_3(),
.F2Adef_R_18_0(),
.F2Adef_R_18_1(),
.F2Adef_R_18_2(),
.F2Adef_R_18_3(),
.F2Adef_R_18_4(),
.F2Adef_R_18_5(),
.F2Adef_R_18_6(),
.F2Adef_R_19_0(),
.F2Adef_R_19_1(),
.F2Adef_R_19_2(),
.F2Adef_R_19_3(),
.F2Adef_R_1_0(),
.F2Adef_R_1_1(),
.F2Adef_R_1_2(),
.F2Adef_R_1_3(),
.F2Adef_R_20_0(),
.F2Adef_R_20_1(),
.F2Adef_R_20_2(),
.F2Adef_R_20_3(),
.F2Adef_R_20_4(),
.F2Adef_R_20_5(),
.F2Adef_R_20_6(),
.F2Adef_R_21_0(),
.F2Adef_R_21_1(),
.F2Adef_R_21_2(),
.F2Adef_R_21_3(),
.F2Adef_R_22_0(),
.F2Adef_R_22_1(),
.F2Adef_R_22_2(),
.F2Adef_R_22_3(),
.F2Adef_R_22_4(),
.F2Adef_R_22_5(),
.F2Adef_R_22_6(),
.F2Adef_R_23_0(),
.F2Adef_R_23_1(),
.F2Adef_R_23_2(),
.F2Adef_R_23_3(),
.F2Adef_R_24_0(),
.F2Adef_R_24_1(),
.F2Adef_R_24_2(),
.F2Adef_R_24_3(),
.F2Adef_R_24_4(),
.F2Adef_R_24_5(),
.F2Adef_R_24_6(),
.F2Adef_R_25_0(),
.F2Adef_R_25_1(),
.F2Adef_R_25_2(),
.F2Adef_R_25_3(),
.F2Adef_R_26_0(),
.F2Adef_R_26_1(),
.F2Adef_R_26_2(),
.F2Adef_R_26_3(),
.F2Adef_R_26_4(),
.F2Adef_R_26_5(),
.F2Adef_R_26_6(),
.F2Adef_R_27_0(),
.F2Adef_R_27_1(),
.F2Adef_R_27_2(),
.F2Adef_R_27_3(),
.F2Adef_R_28_0(),
.F2Adef_R_28_1(),
.F2Adef_R_28_2(),
.F2Adef_R_28_3(),
.F2Adef_R_28_4(),
.F2Adef_R_28_5(),
.F2Adef_R_28_6(),
.F2Adef_R_29_0(),
.F2Adef_R_29_1(),
.F2Adef_R_29_2(),
.F2Adef_R_29_3(),
.F2Adef_R_2_0(),
.F2Adef_R_2_1(),
.F2Adef_R_2_2(),
.F2Adef_R_2_3(),
.F2Adef_R_2_4(),
.F2Adef_R_2_5(),
.F2Adef_R_2_6(),
.F2Adef_R_30_0(),
.F2Adef_R_30_1(),
.F2Adef_R_30_2(),
.F2Adef_R_30_3(),
.F2Adef_R_30_4(),
.F2Adef_R_30_5(),
.F2Adef_R_30_6(),
.F2Adef_R_31_0(),
.F2Adef_R_31_1(),
.F2Adef_R_31_2(),
.F2Adef_R_31_3(),
.F2Adef_R_32_0(),
.F2Adef_R_32_1(),
.F2Adef_R_32_2(),
.F2Adef_R_32_3(),
.F2Adef_R_32_4(),
.F2Adef_R_32_5(),
.F2Adef_R_32_6(),
.F2Adef_R_3_0(),
.F2Adef_R_3_1(),
.F2Adef_R_3_2(),
.F2Adef_R_3_3(),
.F2Adef_R_4_0(),
.F2Adef_R_4_1(),
.F2Adef_R_4_2(),
.F2Adef_R_4_3(),
.F2Adef_R_4_4(),
.F2Adef_R_4_5(),
.F2Adef_R_4_6(),
.F2Adef_R_5_0(),
.F2Adef_R_5_1(),
.F2Adef_R_5_2(),
.F2Adef_R_5_3(),
.F2Adef_R_6_0(),
.F2Adef_R_6_1(),
.F2Adef_R_6_2(),
.F2Adef_R_6_3(),
.F2Adef_R_6_4(),
.F2Adef_R_6_5(),
.F2Adef_R_6_6(),
.F2Adef_R_7_0(),
.F2Adef_R_7_1(),
.F2Adef_R_7_2(),
.F2Adef_R_7_3(),
.F2Adef_R_8_0(),
.F2Adef_R_8_1(),
.F2Adef_R_8_2(),
.F2Adef_R_8_3(),
.F2Adef_R_8_4(),
.F2Adef_R_8_5(),
.F2Adef_R_8_6(),
.F2Adef_R_9_0(),
.F2Adef_R_9_1(),
.F2Adef_R_9_2(),
.F2Adef_R_9_3(),
.F2Adef_T_10_0(),
.F2Adef_T_10_1(),
.F2Adef_T_10_2(),
.F2Adef_T_10_3(),
.F2Adef_T_10_4(),
.F2Adef_T_10_5(),
.F2Adef_T_10_6(),
.F2Adef_T_11_0(),
.F2Adef_T_11_1(),
.F2Adef_T_11_2(),
.F2Adef_T_11_3(),
.F2Adef_T_12_0(),
.F2Adef_T_12_1(),
.F2Adef_T_12_2(),
.F2Adef_T_12_3(),
.F2Adef_T_12_4(),
.F2Adef_T_12_5(),
.F2Adef_T_12_6(),
.F2Adef_T_13_0(),
.F2Adef_T_13_1(),
.F2Adef_T_13_2(),
.F2Adef_T_13_3(),
.F2Adef_T_14_0(),
.F2Adef_T_14_1(),
.F2Adef_T_14_2(),
.F2Adef_T_14_3(),
.F2Adef_T_14_4(),
.F2Adef_T_14_5(),
.F2Adef_T_14_6(),
.F2Adef_T_15_0(),
.F2Adef_T_15_1(),
.F2Adef_T_15_2(),
.F2Adef_T_15_3(),
.F2Adef_T_16_0(),
.F2Adef_T_16_1(),
.F2Adef_T_16_2(),
.F2Adef_T_16_3(),
.F2Adef_T_16_4(),
.F2Adef_T_16_5(),
.F2Adef_T_16_6(),
.F2Adef_T_17_0(),
.F2Adef_T_17_1(),
.F2Adef_T_17_2(),
.F2Adef_T_17_3(),
.F2Adef_T_18_0(),
.F2Adef_T_18_1(),
.F2Adef_T_18_2(),
.F2Adef_T_18_3(),
.F2Adef_T_18_4(),
.F2Adef_T_18_5(),
.F2Adef_T_18_6(),
.F2Adef_T_19_0(),
.F2Adef_T_19_1(),
.F2Adef_T_19_2(),
.F2Adef_T_19_3(),
.F2Adef_T_1_0(),
.F2Adef_T_1_1(),
.F2Adef_T_1_2(),
.F2Adef_T_1_3(),
.F2Adef_T_20_0(),
.F2Adef_T_20_1(),
.F2Adef_T_20_2(),
.F2Adef_T_20_3(),
.F2Adef_T_20_4(),
.F2Adef_T_20_5(),
.F2Adef_T_20_6(),
.F2Adef_T_21_0(),
.F2Adef_T_21_1(),
.F2Adef_T_21_2(),
.F2Adef_T_21_3(),
.F2Adef_T_22_0(),
.F2Adef_T_22_1(MU1_EFPGA_MATHB_TC_defPin),
.F2Adef_T_22_2(MU1_EFPGA_MATHB_OPER_defPin_1_),
.F2Adef_T_22_3(MU1_EFPGA_MATHB_OPER_defPin_0_),
.F2Adef_T_22_4(MU1_EFPGA_MATHB_COEF_defPin_1_),
.F2Adef_T_22_5(MU1_EFPGA_MATHB_COEF_defPin_0_),
.F2Adef_T_22_6(),
.F2Adef_T_23_0(),
.F2Adef_T_23_1(),
.F2Adef_T_23_2(),
.F2Adef_T_23_3(),
.F2Adef_T_24_0(),
.F2Adef_T_24_1(),
.F2Adef_T_24_2(),
.F2Adef_T_24_3(),
.F2Adef_T_24_4(),
.F2Adef_T_24_5(),
.F2Adef_T_24_6(),
.F2Adef_T_25_0(),
.F2Adef_T_25_1(),
.F2Adef_T_25_2(),
.F2Adef_T_25_3(),
.F2Adef_T_26_0(),
.F2Adef_T_26_1(),
.F2Adef_T_26_2(),
.F2Adef_T_26_3(),
.F2Adef_T_26_4(),
.F2Adef_T_26_5(),
.F2Adef_T_26_6(),
.F2Adef_T_27_0(),
.F2Adef_T_27_1(),
.F2Adef_T_27_2(),
.F2Adef_T_27_3(),
.F2Adef_T_28_0(),
.F2Adef_T_28_1(),
.F2Adef_T_28_2(),
.F2Adef_T_28_3(),
.F2Adef_T_28_4(),
.F2Adef_T_28_5(),
.F2Adef_T_28_6(),
.F2Adef_T_29_0(),
.F2Adef_T_29_1(),
.F2Adef_T_29_2(),
.F2Adef_T_29_3(),
.F2Adef_T_2_0(),
.F2Adef_T_2_1(),
.F2Adef_T_2_2(),
.F2Adef_T_2_3(),
.F2Adef_T_2_4(),
.F2Adef_T_2_5(),
.F2Adef_T_2_6(),
.F2Adef_T_30_0(),
.F2Adef_T_30_1(),
.F2Adef_T_30_2(),
.F2Adef_T_30_3(),
.F2Adef_T_30_4(),
.F2Adef_T_30_5(),
.F2Adef_T_30_6(),
.F2Adef_T_31_0(),
.F2Adef_T_31_1(),
.F2Adef_T_31_2(),
.F2Adef_T_31_3(),
.F2Adef_T_32_0(),
.F2Adef_T_32_1(),
.F2Adef_T_32_2(),
.F2Adef_T_32_3(),
.F2Adef_T_32_4(),
.F2Adef_T_32_5(),
.F2Adef_T_32_6(),
.F2Adef_T_3_0(),
.F2Adef_T_3_1(),
.F2Adef_T_3_2(),
.F2Adef_T_3_3(),
.F2Adef_T_4_0(),
.F2Adef_T_4_1(),
.F2Adef_T_4_2(),
.F2Adef_T_4_3(),
.F2Adef_T_4_4(),
.F2Adef_T_4_5(),
.F2Adef_T_4_6(),
.F2Adef_T_5_0(),
.F2Adef_T_5_1(),
.F2Adef_T_5_2(),
.F2Adef_T_5_3(),
.F2Adef_T_6_0(),
.F2Adef_T_6_1(MU0_EFPGA_MATHB_TC_defPin),
.F2Adef_T_6_2(MU0_EFPGA_MATHB_OPER_defPin_1_),
.F2Adef_T_6_3(MU0_EFPGA_MATHB_OPER_defPin_0_),
.F2Adef_T_6_4(MU0_EFPGA_MATHB_COEF_defPin_1_),
.F2Adef_T_6_5(MU0_EFPGA_MATHB_COEF_defPin_0_),
.F2Adef_T_6_6(),
.F2Adef_T_7_0(),
.F2Adef_T_7_1(),
.F2Adef_T_7_2(),
.F2Adef_T_7_3(),
.F2Adef_T_8_0(),
.F2Adef_T_8_1(),
.F2Adef_T_8_2(),
.F2Adef_T_8_3(),
.F2Adef_T_8_4(),
.F2Adef_T_8_5(),
.F2Adef_T_8_6(),
.F2Adef_T_9_0(),
.F2Adef_T_9_1(),
.F2Adef_T_9_2(),
.F2Adef_T_9_3(),
.F2Areg_B_11_0(),
.F2Areg_B_11_1(),
.F2Areg_B_13_0(),
.F2Areg_B_13_1(),
.F2Areg_B_15_0(),
.F2Areg_B_15_1(),
.F2Areg_B_17_0(),
.F2Areg_B_17_1(),
.F2Areg_B_19_0(),
.F2Areg_B_19_1(),
.F2Areg_B_1_0(),
.F2Areg_B_1_1(),
.F2Areg_B_21_0(),
.F2Areg_B_21_1(),
.F2Areg_B_23_0(),
.F2Areg_B_23_1(),
.F2Areg_B_25_0(),
.F2Areg_B_25_1(),
.F2Areg_B_27_0(),
.F2Areg_B_27_1(),
.F2Areg_B_29_0(),
.F2Areg_B_29_1(),
.F2Areg_B_31_0(),
.F2Areg_B_31_1(),
.F2Areg_B_3_0(),
.F2Areg_B_3_1(),
.F2Areg_B_5_0(),
.F2Areg_B_5_1(),
.F2Areg_B_7_0(),
.F2Areg_B_7_1(),
.F2Areg_B_9_0(),
.F2Areg_B_9_1(),
.F2Areg_L_11_0(),
.F2Areg_L_11_1(),
.F2Areg_L_13_0(),
.F2Areg_L_13_1(),
.F2Areg_L_15_0(),
.F2Areg_L_15_1(),
.F2Areg_L_17_0(),
.F2Areg_L_17_1(),
.F2Areg_L_19_0(),
.F2Areg_L_19_1(),
.F2Areg_L_1_0(),
.F2Areg_L_1_1(),
.F2Areg_L_21_0(),
.F2Areg_L_21_1(),
.F2Areg_L_23_0(),
.F2Areg_L_23_1(),
.F2Areg_L_25_0(),
.F2Areg_L_25_1(),
.F2Areg_L_27_0(),
.F2Areg_L_27_1(),
.F2Areg_L_29_0(),
.F2Areg_L_29_1(),
.F2Areg_L_31_0(),
.F2Areg_L_31_1(),
.F2Areg_L_3_0(),
.F2Areg_L_3_1(),
.F2Areg_L_5_0(),
.F2Areg_L_5_1(),
.F2Areg_L_7_0(),
.F2Areg_L_7_1(),
.F2Areg_L_9_0(),
.F2Areg_L_9_1(),
.F2Areg_R_11_0(),
.F2Areg_R_11_1(),
.F2Areg_R_13_0(),
.F2Areg_R_13_1(),
.F2Areg_R_15_0(),
.F2Areg_R_15_1(),
.F2Areg_R_17_0(),
.F2Areg_R_17_1(),
.F2Areg_R_19_0(),
.F2Areg_R_19_1(),
.F2Areg_R_1_0(),
.F2Areg_R_1_1(),
.F2Areg_R_21_0(),
.F2Areg_R_21_1(),
.F2Areg_R_23_0(),
.F2Areg_R_23_1(),
.F2Areg_R_25_0(),
.F2Areg_R_25_1(),
.F2Areg_R_27_0(),
.F2Areg_R_27_1(),
.F2Areg_R_29_0(),
.F2Areg_R_29_1(),
.F2Areg_R_31_0(),
.F2Areg_R_31_1(),
.F2Areg_R_3_0(),
.F2Areg_R_3_1(),
.F2Areg_R_5_0(),
.F2Areg_R_5_1(),
.F2Areg_R_7_0(),
.F2Areg_R_7_1(),
.F2Areg_R_9_0(),
.F2Areg_R_9_1(),
.F2Areg_T_11_0(),
.F2Areg_T_11_1(),
.F2Areg_T_13_0(),
.F2Areg_T_13_1(),
.F2Areg_T_15_0(),
.F2Areg_T_15_1(),
.F2Areg_T_17_0(),
.F2Areg_T_17_1(),
.F2Areg_T_19_0(),
.F2Areg_T_19_1(),
.F2Areg_T_1_0(),
.F2Areg_T_1_1(),
.F2Areg_T_21_0(),
.F2Areg_T_21_1(),
.F2Areg_T_23_0(),
.F2Areg_T_23_1(),
.F2Areg_T_25_0(),
.F2Areg_T_25_1(),
.F2Areg_T_27_0(),
.F2Areg_T_27_1(),
.F2Areg_T_29_0(),
.F2Areg_T_29_1(),
.F2Areg_T_31_0(),
.F2Areg_T_31_1(),
.F2Areg_T_3_0(),
.F2Areg_T_3_1(),
.F2Areg_T_5_0(),
.F2Areg_T_5_1(),
.F2Areg_T_7_0(),
.F2Areg_T_7_1(),
.F2Areg_T_9_0(),
.F2Areg_T_9_1(),
.BL_DOUT_0_(BL_DOUT_0_),
.BL_DOUT_10_(BL_DOUT_10_),
.BL_DOUT_11_(BL_DOUT_11_),
.BL_DOUT_12_(BL_DOUT_12_),
.BL_DOUT_13_(BL_DOUT_13_),
.BL_DOUT_14_(BL_DOUT_14_),
.BL_DOUT_15_(BL_DOUT_15_),
.BL_DOUT_16_(BL_DOUT_16_),
.BL_DOUT_17_(BL_DOUT_17_),
.BL_DOUT_18_(BL_DOUT_18_),
.BL_DOUT_19_(BL_DOUT_19_),
.BL_DOUT_1_(BL_DOUT_1_),
.BL_DOUT_20_(BL_DOUT_20_),
.BL_DOUT_21_(BL_DOUT_21_),
.BL_DOUT_22_(BL_DOUT_22_),
.BL_DOUT_23_(BL_DOUT_23_),
.BL_DOUT_24_(BL_DOUT_24_),
.BL_DOUT_25_(BL_DOUT_25_),
.BL_DOUT_26_(BL_DOUT_26_),
.BL_DOUT_27_(BL_DOUT_27_),
.BL_DOUT_28_(BL_DOUT_28_),
.BL_DOUT_29_(BL_DOUT_29_),
.BL_DOUT_2_(BL_DOUT_2_),
.BL_DOUT_30_(BL_DOUT_30_),
.BL_DOUT_31_(BL_DOUT_31_),
.BL_DOUT_3_(BL_DOUT_3_),
.BL_DOUT_4_(BL_DOUT_4_),
.BL_DOUT_5_(BL_DOUT_5_),
.BL_DOUT_6_(BL_DOUT_6_),
.BL_DOUT_7_(BL_DOUT_7_),
.BL_DOUT_8_(BL_DOUT_8_),
.BL_DOUT_9_(BL_DOUT_9_),
.FB_SPE_OUT_0_(FB_SPE_OUT_0_),
.FB_SPE_OUT_1_(FB_SPE_OUT_1_),
.FB_SPE_OUT_2_(FB_SPE_OUT_2_),
.FB_SPE_OUT_3_(FB_SPE_OUT_3_),
.PARALLEL_CFG(PARALLEL_CFG)
);

endmodule
