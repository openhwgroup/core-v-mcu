module a2_bootrom
 #(
 parameter ADDR_WIDTH=32,
 parameter DATA_WIDTH=32
 )
 (
 input logic 		  CLK,
 input logic 		  CEN,
 input logic [ADDR_WIDTH-1:0]  A,
 output logic [DATA_WIDTH-1:0] Q
 );
 logic [31:0] 		  value;
 assign Q = value;
 always @(posedge CLK) begin
  case (A)
  0: value <= 32'h09C0006F;
  1: value <= 32'h0980006F;
  2: value <= 32'h0940006F;
  3: value <= 32'h0900006F;
  4: value <= 32'h08C0006F;
  5: value <= 32'h0880006F;
  6: value <= 32'h0840006F;
  7: value <= 32'h0800006F;
  8: value <= 32'h07C0006F;
  9: value <= 32'h0780006F;
  10: value <= 32'h0740006F;
  11: value <= 32'h0700006F;
  12: value <= 32'h06C0006F;
  13: value <= 32'h0680006F;
  14: value <= 32'h0640006F;
  15: value <= 32'h0600006F;
  16: value <= 32'h05C0006F;
  17: value <= 32'h0580006F;
  18: value <= 32'h0540006F;
  19: value <= 32'h0500006F;
  20: value <= 32'h04C0006F;
  21: value <= 32'h0480006F;
  22: value <= 32'h0440006F;
  23: value <= 32'h0400006F;
  24: value <= 32'h03C0006F;
  25: value <= 32'h0380006F;
  26: value <= 32'h0340006F;
  27: value <= 32'h0300006F;
  28: value <= 32'h02C0006F;
  29: value <= 32'h0280006F;
  30: value <= 32'h0240006F;
  31: value <= 32'h0200006F;
  32: value <= 32'h0080006F;
  33: value <= 32'h0000006F;
  34: value <= 32'h0207E117;
  35: value <= 32'hFE410113;
  36: value <= 32'h3680006F;
  37: value <= 32'h00060113;
  38: value <= 32'h00058067;
  39: value <= 32'h30200073;
  40: value <= 32'hCA09832A;
  41: value <= 32'h00058383;
  42: value <= 32'h00730023;
  43: value <= 32'h0305167D;
  44: value <= 32'hFA6D0585;
  45: value <= 32'h15F98082;
  46: value <= 32'h114105C2;
  47: value <= 32'hC42281C1;
  48: value <= 32'h842AC606;
  49: value <= 32'h47832A95;
  50: value <= 32'h47030014;
  51: value <= 32'h07A20004;
  52: value <= 32'h67298FD9;
  53: value <= 32'h50770713;
  54: value <= 32'h08E79B63;
  55: value <= 32'h00644783;
  56: value <= 32'h02400713;
  57: value <= 32'h02E79863;
  58: value <= 32'h00344703;
  59: value <= 32'h00244783;
  60: value <= 32'h00544503;
  61: value <= 32'h8F5D0722;
  62: value <= 32'h00444783;
  63: value <= 32'h00744603;
  64: value <= 32'h00840593;
  65: value <= 32'h40B24422;
  66: value <= 32'h8FD907C2;
  67: value <= 32'h8D5D0562;
  68: value <= 32'hB7790141;
  69: value <= 32'h02600713;
  70: value <= 32'h04E79B63;
  71: value <= 32'h1A001537;
  72: value <= 32'h8E850513;
  73: value <= 32'h47032249;
  74: value <= 32'h47830034;
  75: value <= 32'h45030024;
  76: value <= 32'h07220054;
  77: value <= 32'h47838F5D;
  78: value <= 32'h05620044;
  79: value <= 32'h8FD907C2;
  80: value <= 32'h2AC18D5D;
  81: value <= 32'h1A001537;
  82: value <= 32'h92850513;
  83: value <= 32'h47832AA9;
  84: value <= 32'h47030034;
  85: value <= 32'h07A20024;
  86: value <= 32'h47038FD9;
  87: value <= 32'h07420044;
  88: value <= 32'h47838F5D;
  89: value <= 32'h07E20054;
  90: value <= 32'h97828FD9;
  91: value <= 32'h40B2A001;
  92: value <= 32'h01414422;
  93: value <= 32'h11418082;
  94: value <= 32'hC422C606;
  95: value <= 32'hC04AC226;
  96: value <= 32'hC12D240D;
  97: value <= 32'h1C07E7B7;
  98: value <= 32'h84234705;
  99: value <= 32'h2421C6E7;
  100: value <= 32'h02000793;
  101: value <= 32'h00F51A63;
  102: value <= 32'h40B24422;
  103: value <= 32'h49024492;
  104: value <= 32'h02100513;
  105: value <= 32'hA4210141;
  106: value <= 32'h079322FD;
  107: value <= 32'h1B630230;
  108: value <= 32'hE4B702F5;
  109: value <= 32'h44011C07;
  110: value <= 32'h92848913;
  111: value <= 32'h2A75A809;
  112: value <= 32'h008907B3;
  113: value <= 32'h04420405;
  114: value <= 32'h00A78023;
  115: value <= 32'h2A6D8041;
  116: value <= 32'h85A2F57D;
  117: value <= 32'h40B24422;
  118: value <= 32'h85134902;
  119: value <= 32'h44929284;
  120: value <= 32'hBDD10141;
  121: value <= 32'h442240B2;
  122: value <= 32'h49024492;
  123: value <= 32'h80820141;
  124: value <= 32'h1C07E737;
  125: value <= 32'h07136585;
  126: value <= 32'h4601A287;
  127: value <= 32'h02158593;
  128: value <= 32'h10000513;
  129: value <= 32'h00861793;
  130: value <= 32'h83C107C2;
  131: value <= 32'h981346A1;
  132: value <= 32'h58130107;
  133: value <= 32'h07864108;
  134: value <= 32'h00085363;
  135: value <= 32'h16FD8FAD;
  136: value <= 32'hF69307C2;
  137: value <= 32'h83C10FF6;
  138: value <= 32'h1023F2FD;
  139: value <= 32'h060500F7;
  140: value <= 32'h19E30709;
  141: value <= 32'h8082FCA6;
  142: value <= 32'hE63767C1;
  143: value <= 32'h86AA1C07;
  144: value <= 32'h85134701;
  145: value <= 32'h0613FFF7;
  146: value <= 32'h4363A286;
  147: value <= 32'h808200B7;
  148: value <= 32'h00E68833;
  149: value <= 32'h00084803;
  150: value <= 32'h00855793;
  151: value <= 32'hC7B30705;
  152: value <= 32'h07860107;
  153: value <= 32'hD80397B2;
  154: value <= 32'h17930007;
  155: value <= 32'h07C20085;
  156: value <= 32'h453383C1;
  157: value <= 32'hBFD100F8;
  158: value <= 32'hC62A1101;
  159: value <= 32'h45850070;
  160: value <= 32'hCE064505;
  161: value <= 32'h40F22535;
  162: value <= 32'h80826105;
  163: value <= 32'h45351141;
  164: value <= 32'h37DDC606;
  165: value <= 32'h452940B2;
  166: value <= 32'hBFF90141;
  167: value <= 32'h136347A9;
  168: value <= 32'hB7ED00F5;
  169: value <= 32'h1141BFD1;
  170: value <= 32'hC606C422;
  171: value <= 32'h0503842A;
  172: value <= 32'hE5090004;
  173: value <= 32'h442240B2;
  174: value <= 32'h80820141;
  175: value <= 32'h040537C5;
  176: value <= 32'h5793B7FD;
  177: value <= 32'h11410045;
  178: value <= 32'hC4228BBD;
  179: value <= 32'h842AC606;
  180: value <= 32'h03900713;
  181: value <= 32'h03078513;
  182: value <= 32'h00A75463;
  183: value <= 32'h05778513;
  184: value <= 32'h883D3F75;
  185: value <= 32'h03040513;
  186: value <= 32'h03900793;
  187: value <= 32'h00A7D463;
  188: value <= 32'h05740513;
  189: value <= 32'h40B24422;
  190: value <= 32'hB74D0141;
  191: value <= 32'hC4221141;
  192: value <= 32'h8121842A;
  193: value <= 32'h3F75C606;
  194: value <= 32'h44228522;
  195: value <= 32'h014140B2;
  196: value <= 32'h1141BF4D;
  197: value <= 32'h842AC422;
  198: value <= 32'hC6068141;
  199: value <= 32'h852237C5;
  200: value <= 32'h40B24422;
  201: value <= 32'hBFD90141;
  202: value <= 32'h1A1077B7;
  203: value <= 32'h75134388;
  204: value <= 32'h808207F5;
  205: value <= 32'h1A107737;
  206: value <= 32'h00074783;
  207: value <= 32'h07F57513;
  208: value <= 32'hF807F793;
  209: value <= 32'h00238FC9;
  210: value <= 32'h808200F7;
  211: value <= 32'h1F634785;
  212: value <= 32'h773700F5;
  213: value <= 32'h47831A10;
  214: value <= 32'hE7930047;
  215: value <= 32'h02230017;
  216: value <= 32'h77B700F7;
  217: value <= 32'h43C81A10;
  218: value <= 32'h80828905;
  219: value <= 32'h7737F97D;
  220: value <= 32'h47831A10;
  221: value <= 32'h9BF90047;
  222: value <= 32'h77B7B7DD;
  223: value <= 32'hA5031A10;
  224: value <= 32'h75130847;
  225: value <= 32'h80820FF5;
  226: value <= 32'h1A1077B7;
  227: value <= 32'h0907A503;
  228: value <= 32'h0FF57513;
  229: value <= 32'h77B78082;
  230: value <= 32'h43A81A10;
  231: value <= 32'h0FF57513;
  232: value <= 32'h77B78082;
  233: value <= 32'h43E81A10;
  234: value <= 32'h0FF57513;
  235: value <= 32'h77B78082;
  236: value <= 32'hC7A81A10;
  237: value <= 32'hD5B78082;
  238: value <= 32'h11411C07;
  239: value <= 32'h85934641;
  240: value <= 32'h45014085;
  241: value <= 32'h2EF1C606;
  242: value <= 32'h1C07D7B7;
  243: value <= 32'h40C7A603;
  244: value <= 32'hCE6347BD;
  245: value <= 32'hCE1100C7;
  246: value <= 32'h061240B2;
  247: value <= 32'hD5B70642;
  248: value <= 32'h82411C07;
  249: value <= 32'h41858593;
  250: value <= 32'h01414541;
  251: value <= 32'h4641AE5D;
  252: value <= 32'h40B2B7E5;
  253: value <= 32'h80820141;
  254: value <= 32'h1C0107B7;
  255: value <= 32'h715D439C;
  256: value <= 32'h1A1047B7;
  257: value <= 32'hC6864505;
  258: value <= 32'hC2A6C4A2;
  259: value <= 32'h0C47A403;
  260: value <= 32'hDE4EC0CA;
  261: value <= 32'hDA56DC52;
  262: value <= 32'hD65ED85A;
  263: value <= 32'hD266D462;
  264: value <= 32'hCE6ED06A;
  265: value <= 32'h37093725;
  266: value <= 32'h06200793;
  267: value <= 32'h05638805;
  268: value <= 32'h051300F5;
  269: value <= 32'h3DFD0620;
  270: value <= 32'h859365F1;
  271: value <= 32'h45052005;
  272: value <= 32'h15372131;
  273: value <= 32'h05131A00;
  274: value <= 32'h3DB18F85;
  275: value <= 32'h0E040163;
  276: value <= 32'h1A001537;
  277: value <= 32'h91050513;
  278: value <= 32'h25B735B9;
  279: value <= 32'h85930026;
  280: value <= 32'h45015A05;
  281: value <= 32'h45812A4D;
  282: value <= 32'h2C854501;
  283: value <= 32'h45014581;
  284: value <= 32'h002824F9;
  285: value <= 32'hE4092AE9;
  286: value <= 32'h02E00793;
  287: value <= 32'h00F10423;
  288: value <= 32'h000104A3;
  289: value <= 32'h14040D63;
  290: value <= 32'h1C07C9B7;
  291: value <= 32'h84136785;
  292: value <= 32'h64890009;
  293: value <= 32'h00940933;
  294: value <= 32'h2023943E;
  295: value <= 32'h2E2392F9;
  296: value <= 32'h22239009;
  297: value <= 32'h22239209;
  298: value <= 32'h37314004;
  299: value <= 32'h92092783;
  300: value <= 32'h40C42803;
  301: value <= 32'h1C07D6B7;
  302: value <= 32'h1C07EA37;
  303: value <= 32'h1C07D937;
  304: value <= 32'hFFF78893;
  305: value <= 32'h40F00633;
  306: value <= 32'h42068693;
  307: value <= 32'h07B74581;
  308: value <= 32'h0A131C00;
  309: value <= 32'h0913000A;
  310: value <= 32'h84930009;
  311: value <= 32'h9D639284;
  312: value <= 32'h67090505;
  313: value <= 32'h670597BA;
  314: value <= 32'h9007AE23;
  315: value <= 32'h9207A223;
  316: value <= 32'h92E7A023;
  317: value <= 32'h1C07D437;
  318: value <= 32'h04133D7D;
  319: value <= 32'h4A814184;
  320: value <= 32'h01000CB7;
  321: value <= 32'h40C92783;
  322: value <= 32'h04FAED63;
  323: value <= 32'h1A001537;
  324: value <= 32'h92C50513;
  325: value <= 32'h25033B49;
  326: value <= 32'h3BE54109;
  327: value <= 32'h1A001537;
  328: value <= 32'h92850513;
  329: value <= 32'h27833349;
  330: value <= 32'h97824109;
  331: value <= 32'h1537A001;
  332: value <= 32'h05131A00;
  333: value <= 32'hB70D9145;
  334: value <= 32'hFFC6A703;
  335: value <= 32'h00E7E963;
  336: value <= 32'h953A4288;
  337: value <= 32'h00A7E963;
  338: value <= 32'h06C10585;
  339: value <= 32'h8533BF49;
  340: value <= 32'h7BE30097;
  341: value <= 32'h429CFEA7;
  342: value <= 32'h9746973E;
  343: value <= 32'h00C777B3;
  344: value <= 32'h17B7B7E5;
  345: value <= 32'h85131A00;
  346: value <= 32'h3B359187;
  347: value <= 32'h33558556;
  348: value <= 32'h1A0017B7;
  349: value <= 32'h93478513;
  350: value <= 32'h4048333D;
  351: value <= 32'h3B514B01;
  352: value <= 32'h00442D83;
  353: value <= 32'h00042C03;
  354: value <= 32'h00842B83;
  355: value <= 32'hE40007B7;
  356: value <= 32'h00FD8D33;
  357: value <= 32'h65634450;
  358: value <= 32'h0A8500CB;
  359: value <= 32'hB79D0441;
  360: value <= 32'h920A2483;
  361: value <= 32'h009BF563;
  362: value <= 32'h003B8493;
  363: value <= 32'h961398F1;
  364: value <= 32'h82410104;
  365: value <= 32'h019D7B63;
  366: value <= 32'h856285EE;
  367: value <= 32'h9DA622DD;
  368: value <= 32'h8BB39C26;
  369: value <= 32'h0B05409B;
  370: value <= 32'h8593B7F1;
  371: value <= 32'h85620009;
  372: value <= 32'h86262AC9;
  373: value <= 32'h00098593;
  374: value <= 32'h34D9856E;
  375: value <= 32'h3909B7CD;
  376: value <= 32'h1A1047B7;
  377: value <= 32'hDBF84705;
  378: value <= 32'h0007A937;
  379: value <= 32'h1A1044B7;
  380: value <= 32'hEA374985;
  381: value <= 32'h04131C07;
  382: value <= 32'h58FC1209;
  383: value <= 32'h01378463;
  384: value <= 32'h3B0158E8;
  385: value <= 32'h3E85147D;
  386: value <= 32'h4783F86D;
  387: value <= 32'hF7E5C68A;
  388: value <= 32'h39510028;
  389: value <= 32'h2737B7CD;
  390: value <= 32'h47141A10;
  391: value <= 32'h95334791;
  392: value <= 32'h8EC900A7;
  393: value <= 32'h4714C714;
  394: value <= 32'hFFF54793;
  395: value <= 32'hC71C8FF5;
  396: value <= 32'h8D5D431C;
  397: value <= 32'h004C57B7;
  398: value <= 32'hB4078793;
  399: value <= 32'h02B7D7B3;
  400: value <= 32'hE737C308;
  401: value <= 32'h45011C07;
  402: value <= 32'hC6F704A3;
  403: value <= 32'h26378082;
  404: value <= 32'h47031A10;
  405: value <= 32'hE6B71886;
  406: value <= 32'h07931C07;
  407: value <= 32'h9B3D1806;
  408: value <= 32'h18E60423;
  409: value <= 32'h19864703;
  410: value <= 32'h0C239B3D;
  411: value <= 32'h470318E6;
  412: value <= 32'h9B3D1A86;
  413: value <= 32'h1AE60423;
  414: value <= 32'hC696C683;
  415: value <= 32'h1C07E737;
  416: value <= 32'hC2870713;
  417: value <= 32'h06B7C314;
  418: value <= 32'hC3541000;
  419: value <= 32'h200706B7;
  420: value <= 32'h09F68693;
  421: value <= 32'h06B7C714;
  422: value <= 32'h068D7047;
  423: value <= 32'h06B7C754;
  424: value <= 32'h06859000;
  425: value <= 32'h2023CB14;
  426: value <= 32'h469118A6;
  427: value <= 32'h4683C3D4;
  428: value <= 32'hE6931886;
  429: value <= 32'h04230106;
  430: value <= 32'hD39818D6;
  431: value <= 32'hD3D84751;
  432: value <= 32'h1A864703;
  433: value <= 32'h01076713;
  434: value <= 32'h1AE60423;
  435: value <= 32'h1A102737;
  436: value <= 32'h18070793;
  437: value <= 32'hFFED43DC;
  438: value <= 32'h27B78082;
  439: value <= 32'h87930034;
  440: value <= 32'h953E0437;
  441: value <= 32'h4783051E;
  442: value <= 32'hE7370285;
  443: value <= 32'h47031C07;
  444: value <= 32'h9BBDC697;
  445: value <= 32'h02F50423;
  446: value <= 32'h02854783;
  447: value <= 32'h0407E793;
  448: value <= 32'h02F50423;
  449: value <= 32'h1C07E7B7;
  450: value <= 32'hC2878793;
  451: value <= 32'h0737C398;
  452: value <= 32'h8DD91000;
  453: value <= 32'h20070737;
  454: value <= 32'h06670713;
  455: value <= 32'h0737C798;
  456: value <= 32'h07059000;
  457: value <= 32'hC3CCD11C;
  458: value <= 32'h47C1C7D8;
  459: value <= 32'h4783D15C;
  460: value <= 32'hE7930285;
  461: value <= 32'h04230107;
  462: value <= 32'h450102F5;
  463: value <= 32'h27B78082;
  464: value <= 32'h87930034;
  465: value <= 32'h953E0437;
  466: value <= 32'h4783051E;
  467: value <= 32'hE7370285;
  468: value <= 32'h47031C07;
  469: value <= 32'h9BBDC697;
  470: value <= 32'h02F50423;
  471: value <= 32'h02854783;
  472: value <= 32'h0407E793;
  473: value <= 32'h02F50423;
  474: value <= 32'h1C07E7B7;
  475: value <= 32'hC2878793;
  476: value <= 32'h0737C398;
  477: value <= 32'h8DD91000;
  478: value <= 32'h20070737;
  479: value <= 32'h09970713;
  480: value <= 32'h0737C798;
  481: value <= 32'h07059000;
  482: value <= 32'hC3CCD11C;
  483: value <= 32'h47C1C7D8;
  484: value <= 32'h4783D15C;
  485: value <= 32'hE7930285;
  486: value <= 32'h04230107;
  487: value <= 32'h450102F5;
  488: value <= 32'h28378082;
  489: value <= 32'h47031A10;
  490: value <= 32'hE6B71888;
  491: value <= 32'h08B71C07;
  492: value <= 32'h9B3D2007;
  493: value <= 32'h18E80423;
  494: value <= 32'h19884703;
  495: value <= 32'h200F0337;
  496: value <= 32'h18080793;
  497: value <= 32'h0C239B3D;
  498: value <= 32'h470318E8;
  499: value <= 32'h9B3D1A88;
  500: value <= 32'h1AE80423;
  501: value <= 32'hC696C683;
  502: value <= 32'h1C07E737;
  503: value <= 32'hC2870713;
  504: value <= 32'h06B7C314;
  505: value <= 32'hC3541000;
  506: value <= 32'h00388693;
  507: value <= 32'h5693C714;
  508: value <= 32'h06C20085;
  509: value <= 32'h751382C1;
  510: value <= 32'hE6B30FF5;
  511: value <= 32'h65330066;
  512: value <= 32'hC7540115;
  513: value <= 32'h0693CB08;
  514: value <= 32'h0537FFF6;
  515: value <= 32'h8EC97047;
  516: value <= 32'h06B7CB54;
  517: value <= 32'h06859000;
  518: value <= 32'h2023CF14;
  519: value <= 32'hC3D018B8;
  520: value <= 32'h18884683;
  521: value <= 32'h0106E693;
  522: value <= 32'h18D80423;
  523: value <= 32'h4771D398;
  524: value <= 32'h4703D3D8;
  525: value <= 32'h67131A88;
  526: value <= 32'h04230107;
  527: value <= 32'h27371AE8;
  528: value <= 32'h07931A10;
  529: value <= 32'h43DC1807;
  530: value <= 32'h8082FFED;
  531: value <= 32'h1A102737;
  532: value <= 32'h47854714;
  533: value <= 32'h00A797B3;
  534: value <= 32'hC7148EDD;
  535: value <= 32'hC6934710;
  536: value <= 32'h8EF1FFF7;
  537: value <= 32'h4314C714;
  538: value <= 32'hC31C8FD5;
  539: value <= 32'h003427B7;
  540: value <= 32'h04178793;
  541: value <= 32'h57B7953E;
  542: value <= 32'h8793004C;
  543: value <= 32'hD7B3B407;
  544: value <= 32'h051E02B7;
  545: value <= 32'h83C107C2;
  546: value <= 32'h02F51323;
  547: value <= 32'hE793515C;
  548: value <= 32'hD15C0067;
  549: value <= 32'hE793515C;
  550: value <= 32'hD15C0107;
  551: value <= 32'hE793515C;
  552: value <= 32'hD15C1007;
  553: value <= 32'hE793515C;
  554: value <= 32'hD15C2007;
  555: value <= 32'h80824501;
  556: value <= 32'h003427B7;
  557: value <= 32'h04178793;
  558: value <= 32'h1793953E;
  559: value <= 32'h45010075;
  560: value <= 32'hEF114BD8;
  561: value <= 32'hCBCCCB90;
  562: value <= 32'h0187C703;
  563: value <= 32'h01076713;
  564: value <= 32'h00E78C23;
  565: value <= 32'hE7114BD8;
  566: value <= 32'h81410542;
  567: value <= 32'h05058082;
  568: value <= 32'h0505B7C5;
  569: value <= 32'h0000BFC5;
  570: value <= 32'h4332490A;
  571: value <= 32'h204C4220;
  572: value <= 32'h20504D4A;
  573: value <= 32'h00000000;
  574: value <= 32'h2032410A;
  575: value <= 32'h746F6F42;
  576: value <= 32'h64616F6C;
  577: value <= 32'h42207265;
  578: value <= 32'h73746F6F;
  579: value <= 32'h003D6C65;
  580: value <= 32'h00000031;
  581: value <= 32'h00000030;
  582: value <= 32'h616F4C0A;
  583: value <= 32'h676E6964;
  584: value <= 32'h63655320;
  585: value <= 32'h6E6F6974;
  586: value <= 32'h00000020;
  587: value <= 32'h6D754A0A;
  588: value <= 32'h676E6970;
  589: value <= 32'h206F7420;
  590: value <= 32'h00000000;
  default: value <= 0;
   endcase
  end
endmodule    
