`define INFO                      'h0000
`define JTAGREG                   'h0074
`define CORESTATUS                'h00A0
`define CS_RO                     'h00C0
`define BOOTSEL                   'h00C4
`define CLKSEL                    'h00C8
`define CLK_DIV_CLU               'h00D8
`define SEL_CLK_DC_FIFO_EFPGA     'h00E0
`define CLK_GATING_DC_FIFO_EFPGA  'h00E4
`define RESET_TYPE1_EFPGA         'h00E8
`define ENABLE_IN_OUT_EFPGA       'h00EC
`define IO_CTRL                   'h0400
