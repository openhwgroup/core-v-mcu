//{{{
wire                    MU0_EFPGA2MATHB_CLK;    // From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire                    MU0_EFPGA_MATHB_CLK_EN; // From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [31:0]             MU0_EFPGA_MATHB_COEF_DATA;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU0_EFPGA_MATHB_COEF_SEL;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [1:0]              MU0_EFPGA_MATHB_COEF_defPin;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire [1:0]              MU0_EFPGA_MATHB_DATAOUT_SEL;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU0_EFPGA_MATHB_MAC_ACC_CLEAR;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire                    MU0_EFPGA_MATHB_MAC_ACC_RND;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire                    MU0_EFPGA_MATHB_MAC_ACC_SAT;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [5:0]              MU0_EFPGA_MATHB_MAC_OUT_SEL;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire [31:0]             MU0_EFPGA_MATHB_OPER_DATA;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU0_EFPGA_MATHB_OPER_SEL;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [1:0]              MU0_EFPGA_MATHB_OPER_defPin;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU0_EFPGA_MATHB_TC_defPin;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire                    MU0_EFPGA_TPRAM_COEF_POWERDN;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [11:0]             MU0_EFPGA_TPRAM_COEF_R_ADDR;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU0_EFPGA_TPRAM_COEF_R_CLK;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [1:0]              MU0_EFPGA_TPRAM_COEF_R_MODE;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU0_EFPGA_TPRAM_COEF_WDSEL;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire                    MU0_EFPGA_TPRAM_COEF_WE;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [11:0]             MU0_EFPGA_TPRAM_COEF_W_ADDR;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU0_EFPGA_TPRAM_COEF_W_CLK;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [31:0]             MU0_EFPGA_TPRAM_COEF_W_DATA;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire [1:0]              MU0_EFPGA_TPRAM_COEF_W_MODE;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU0_EFPGA_TPRAM_OPER_POWERDN;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [11:0]             MU0_EFPGA_TPRAM_OPER_R_ADDR;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU0_EFPGA_TPRAM_OPER_R_CLK;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [1:0]              MU0_EFPGA_TPRAM_OPER_R_MODE;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU0_EFPGA_TPRAM_OPER_WDSEL;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire                    MU0_EFPGA_TPRAM_OPER_WE;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [11:0]             MU0_EFPGA_TPRAM_OPER_W_ADDR;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU0_EFPGA_TPRAM_OPER_W_CLK;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [31:0]             MU0_EFPGA_TPRAM_OPER_W_DATA;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire [1:0]              MU0_EFPGA_TPRAM_OPER_W_MODE;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire [31:0]             MU0_MATHB_EFPGA_MAC_OUT;// From U0_MATH_UNIT of MATH_UNIT.v
wire [31:0]             MU0_TPRAM_EFPGA_COEF_R_DATA;// From U0_MATH_UNIT of MATH_UNIT.v
wire [31:0]             MU0_TPRAM_EFPGA_OPER_R_DATA;// From U0_MATH_UNIT of MATH_UNIT.v
wire                    MU1_EFPGA2MATHB_CLK;    // From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire                    MU1_EFPGA_MATHB_CLK_EN; // From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [31:0]             MU1_EFPGA_MATHB_COEF_DATA;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU1_EFPGA_MATHB_COEF_SEL;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [1:0]              MU1_EFPGA_MATHB_COEF_defPin;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire [1:0]              MU1_EFPGA_MATHB_DATAOUT_SEL;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU1_EFPGA_MATHB_MAC_ACC_CLEAR;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire                    MU1_EFPGA_MATHB_MAC_ACC_RND;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire                    MU1_EFPGA_MATHB_MAC_ACC_SAT;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [5:0]              MU1_EFPGA_MATHB_MAC_OUT_SEL;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire [31:0]             MU1_EFPGA_MATHB_OPER_DATA;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU1_EFPGA_MATHB_OPER_SEL;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [1:0]              MU1_EFPGA_MATHB_OPER_defPin;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU1_EFPGA_MATHB_TC_defPin;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire                    MU1_EFPGA_TPRAM_COEF_POWERDN;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [11:0]             MU1_EFPGA_TPRAM_COEF_R_ADDR;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU1_EFPGA_TPRAM_COEF_R_CLK;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [1:0]              MU1_EFPGA_TPRAM_COEF_R_MODE;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU1_EFPGA_TPRAM_COEF_WDSEL;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire                    MU1_EFPGA_TPRAM_COEF_WE;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [11:0]             MU1_EFPGA_TPRAM_COEF_W_ADDR;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU1_EFPGA_TPRAM_COEF_W_CLK;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [31:0]             MU1_EFPGA_TPRAM_COEF_W_DATA;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire [1:0]              MU1_EFPGA_TPRAM_COEF_W_MODE;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU1_EFPGA_TPRAM_OPER_POWERDN;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [11:0]             MU1_EFPGA_TPRAM_OPER_R_ADDR;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU1_EFPGA_TPRAM_OPER_R_CLK;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [1:0]              MU1_EFPGA_TPRAM_OPER_R_MODE;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU1_EFPGA_TPRAM_OPER_WDSEL;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire                    MU1_EFPGA_TPRAM_OPER_WE;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [11:0]             MU1_EFPGA_TPRAM_OPER_W_ADDR;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire                    MU1_EFPGA_TPRAM_OPER_W_CLK;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v
wire [31:0]             MU1_EFPGA_TPRAM_OPER_W_DATA;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire [1:0]              MU1_EFPGA_TPRAM_OPER_W_MODE;// From U_EFPGA_TOP of QL_eFPGA_ArcticPro2_32X32_GF_22_ETH_ARNOLD_Design.v, ...
wire [31:0]             MU1_MATHB_EFPGA_MAC_OUT;// From U1_MATH_UNIT of MATH_UNIT.v
wire [31:0]             MU1_TPRAM_EFPGA_COEF_R_DATA;// From U1_MATH_UNIT of MATH_UNIT.v
wire [31:0]             MU1_TPRAM_EFPGA_OPER_R_DATA;// From U1_MATH_UNIT of MATH_UNIT.v
//}}}