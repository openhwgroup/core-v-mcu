module a2_bootrom
 #(
 parameter ADDR_WIDTH=32,
 parameter DATA_WIDTH=32
 )
 (
 input logic 		  CLK,
 input logic 		  CEN,
 input logic [ADDR_WIDTH-1:0]  A,
 output logic [DATA_WIDTH-1:0] Q
 );
 logic [31:0] 		  value;
 assign Q = value;
 always @(posedge CLK) begin
  case (A)
  0: value <= 32'h09C0006F;
  1: value <= 32'h0980006F;
  2: value <= 32'h0940006F;
  3: value <= 32'h0900006F;
  4: value <= 32'h08C0006F;
  5: value <= 32'h0880006F;
  6: value <= 32'h0840006F;
  7: value <= 32'h0800006F;
  8: value <= 32'h07C0006F;
  9: value <= 32'h0780006F;
  10: value <= 32'h0740006F;
  11: value <= 32'h0700006F;
  12: value <= 32'h06C0006F;
  13: value <= 32'h0680006F;
  14: value <= 32'h0640006F;
  15: value <= 32'h0600006F;
  16: value <= 32'h05C0006F;
  17: value <= 32'h0580006F;
  18: value <= 32'h0540006F;
  19: value <= 32'h0500006F;
  20: value <= 32'h04C0006F;
  21: value <= 32'h0480006F;
  22: value <= 32'h0440006F;
  23: value <= 32'h0400006F;
  24: value <= 32'h03C0006F;
  25: value <= 32'h0380006F;
  26: value <= 32'h0340006F;
  27: value <= 32'h0300006F;
  28: value <= 32'h02C0006F;
  29: value <= 32'h0280006F;
  30: value <= 32'h0240006F;
  31: value <= 32'h0200006F;
  32: value <= 32'h0080006F;
  33: value <= 32'h0000006F;
  34: value <= 32'h0207E117;
  35: value <= 32'hFE410113;
  36: value <= 32'h5C60006F;
  37: value <= 32'h00060113;
  38: value <= 32'h00058067;
  39: value <= 32'h30200073;
  40: value <= 32'hCA09832A;
  41: value <= 32'h00058383;
  42: value <= 32'h00730023;
  43: value <= 32'h0305167D;
  44: value <= 32'hFA6D0585;
  45: value <= 32'h11018082;
  46: value <= 32'hE937C84A;
  47: value <= 32'hC4521C07;
  48: value <= 32'hC6990A13;
  49: value <= 32'h4983C64E;
  50: value <= 32'hCC22000A;
  51: value <= 32'hCA26CE06;
  52: value <= 32'h842A4785;
  53: value <= 32'hC6990913;
  54: value <= 32'h06F98563;
  55: value <= 32'h00144783;
  56: value <= 32'h00044703;
  57: value <= 32'h8FD907A2;
  58: value <= 32'h07136729;
  59: value <= 32'h92635077;
  60: value <= 32'h478304E7;
  61: value <= 32'h07130064;
  62: value <= 32'h92630240;
  63: value <= 32'h470308E7;
  64: value <= 32'h47830034;
  65: value <= 32'h45030024;
  66: value <= 32'h07220054;
  67: value <= 32'h47838F5D;
  68: value <= 32'h46030044;
  69: value <= 32'h05620074;
  70: value <= 32'h8FD907C2;
  71: value <= 32'h00840593;
  72: value <= 32'h3FBD8D5D;
  73: value <= 32'h00094703;
  74: value <= 32'h05134785;
  75: value <= 32'h00630310;
  76: value <= 32'h40F204F7;
  77: value <= 32'h44D24462;
  78: value <= 32'h49B24942;
  79: value <= 32'h61054A22;
  80: value <= 32'h84AE8082;
  81: value <= 32'h05C215F9;
  82: value <= 32'h22AD81C1;
  83: value <= 32'hC70394A2;
  84: value <= 32'hC783FFE4;
  85: value <= 32'h0722FFF4;
  86: value <= 32'h07C28FD9;
  87: value <= 32'h8FE383C1;
  88: value <= 32'h4783F6A7;
  89: value <= 32'h96E3000A;
  90: value <= 32'h0513FD37;
  91: value <= 32'h44620300;
  92: value <= 32'h44D240F2;
  93: value <= 32'h49B24942;
  94: value <= 32'h61054A22;
  95: value <= 32'h0713AC45;
  96: value <= 32'h91E30260;
  97: value <= 32'h1537FAE7;
  98: value <= 32'h05131A00;
  99: value <= 32'h2A59AF85;
  100: value <= 32'h00344703;
  101: value <= 32'h00244783;
  102: value <= 32'h00544503;
  103: value <= 32'h8F5D0722;
  104: value <= 32'h00444783;
  105: value <= 32'h07C20562;
  106: value <= 32'h8D5D8FD9;
  107: value <= 32'h153722D5;
  108: value <= 32'h05131A00;
  109: value <= 32'h22BDB185;
  110: value <= 32'h00344783;
  111: value <= 32'h00244703;
  112: value <= 32'h8FD907A2;
  113: value <= 32'h00444703;
  114: value <= 32'h8F5D0742;
  115: value <= 32'h00544783;
  116: value <= 32'h8FD907E2;
  117: value <= 32'hA0019782;
  118: value <= 32'hC6061141;
  119: value <= 32'hC226C422;
  120: value <= 32'h2C3DC04A;
  121: value <= 32'hE7B7CD35;
  122: value <= 32'h44051C07;
  123: value <= 32'hC6878423;
  124: value <= 32'h47E52415;
  125: value <= 32'h00F51E63;
  126: value <= 32'h1C07E7B7;
  127: value <= 32'hC60784A3;
  128: value <= 32'h40B24422;
  129: value <= 32'h49024492;
  130: value <= 32'h02100513;
  131: value <= 32'hAC390141;
  132: value <= 32'h07932411;
  133: value <= 32'h17630200;
  134: value <= 32'hE7B700F5;
  135: value <= 32'h84A31C07;
  136: value <= 32'hBFF9C687;
  137: value <= 32'h07932AC5;
  138: value <= 32'h1B630230;
  139: value <= 32'hE4B702F5;
  140: value <= 32'h44011C07;
  141: value <= 32'h92848913;
  142: value <= 32'h2A7DA809;
  143: value <= 32'h008907B3;
  144: value <= 32'h04420405;
  145: value <= 32'h00A78023;
  146: value <= 32'h2A758041;
  147: value <= 32'h85A2F57D;
  148: value <= 32'h40B24422;
  149: value <= 32'h85134902;
  150: value <= 32'h44929284;
  151: value <= 32'hBDA10141;
  152: value <= 32'h442240B2;
  153: value <= 32'h49024492;
  154: value <= 32'h80820141;
  155: value <= 32'h1C07E737;
  156: value <= 32'h07136585;
  157: value <= 32'h4601A287;
  158: value <= 32'h02158593;
  159: value <= 32'h10000513;
  160: value <= 32'h00861793;
  161: value <= 32'h83C107C2;
  162: value <= 32'h981346A1;
  163: value <= 32'h58130107;
  164: value <= 32'h07864108;
  165: value <= 32'h00085363;
  166: value <= 32'h16FD8FAD;
  167: value <= 32'hF69307C2;
  168: value <= 32'h83C10FF6;
  169: value <= 32'h1023F2FD;
  170: value <= 32'h060500F7;
  171: value <= 32'h19E30709;
  172: value <= 32'h8082FCA6;
  173: value <= 32'hE63767C1;
  174: value <= 32'h86AA1C07;
  175: value <= 32'h85134701;
  176: value <= 32'h0613FFF7;
  177: value <= 32'h4363A286;
  178: value <= 32'h808200B7;
  179: value <= 32'h00E68833;
  180: value <= 32'h00084803;
  181: value <= 32'h00855793;
  182: value <= 32'hC7B30705;
  183: value <= 32'h07860107;
  184: value <= 32'hD80397B2;
  185: value <= 32'h17930007;
  186: value <= 32'h07C20085;
  187: value <= 32'h453383C1;
  188: value <= 32'hBFD100F8;
  189: value <= 32'hC62A1101;
  190: value <= 32'h45850070;
  191: value <= 32'hCE064505;
  192: value <= 32'h7C2000EF;
  193: value <= 32'h610540F2;
  194: value <= 32'h11418082;
  195: value <= 32'hC6064535;
  196: value <= 32'h40B237D5;
  197: value <= 32'h01414529;
  198: value <= 32'h47A9BFF1;
  199: value <= 32'h00F51363;
  200: value <= 32'hBFC9B7ED;
  201: value <= 32'hC4221141;
  202: value <= 32'h842AC606;
  203: value <= 32'h00040503;
  204: value <= 32'h40B2E509;
  205: value <= 32'h01414422;
  206: value <= 32'h37C58082;
  207: value <= 32'hB7FD0405;
  208: value <= 32'h00455793;
  209: value <= 32'h8BBD1141;
  210: value <= 32'hC606C422;
  211: value <= 32'h0713842A;
  212: value <= 32'h85130390;
  213: value <= 32'h54630307;
  214: value <= 32'h851300A7;
  215: value <= 32'h3F750577;
  216: value <= 32'h0513883D;
  217: value <= 32'h07930304;
  218: value <= 32'hD4630390;
  219: value <= 32'h051300A7;
  220: value <= 32'h44220574;
  221: value <= 32'h014140B2;
  222: value <= 32'h1141B74D;
  223: value <= 32'h842AC422;
  224: value <= 32'hC6068121;
  225: value <= 32'h85223F75;
  226: value <= 32'h40B24422;
  227: value <= 32'hBF4D0141;
  228: value <= 32'hC4221141;
  229: value <= 32'h8141842A;
  230: value <= 32'h37C5C606;
  231: value <= 32'h44228522;
  232: value <= 32'h014140B2;
  233: value <= 32'h77B7BFD9;
  234: value <= 32'h43881A10;
  235: value <= 32'h07F57513;
  236: value <= 32'h77378082;
  237: value <= 32'h47831A10;
  238: value <= 32'h75130007;
  239: value <= 32'hF79307F5;
  240: value <= 32'h8FC9F807;
  241: value <= 32'h00F70023;
  242: value <= 32'h47858082;
  243: value <= 32'h00F51F63;
  244: value <= 32'h1A107737;
  245: value <= 32'h00474783;
  246: value <= 32'h0017E793;
  247: value <= 32'h00F70223;
  248: value <= 32'h1A1077B7;
  249: value <= 32'h890543C8;
  250: value <= 32'hF97D8082;
  251: value <= 32'h1A107737;
  252: value <= 32'h00474783;
  253: value <= 32'hB7DD9BF9;
  254: value <= 32'h1A1077B7;
  255: value <= 32'h0847A503;
  256: value <= 32'h0FF57513;
  257: value <= 32'h77B78082;
  258: value <= 32'hA5031A10;
  259: value <= 32'h75130907;
  260: value <= 32'h80820FF5;
  261: value <= 32'h1A1077B7;
  262: value <= 32'h751343A8;
  263: value <= 32'h80820FF5;
  264: value <= 32'h1A1077B7;
  265: value <= 32'h751343E8;
  266: value <= 32'h80820FF5;
  267: value <= 32'h1A1077B7;
  268: value <= 32'h8082C7A8;
  269: value <= 32'hC2261141;
  270: value <= 32'h85936485;
  271: value <= 32'hC4224084;
  272: value <= 32'h842A4641;
  273: value <= 32'h450195AA;
  274: value <= 32'h94A2C606;
  275: value <= 32'hA60323A5;
  276: value <= 32'h47BD40C4;
  277: value <= 32'h00C7CE63;
  278: value <= 32'h6585CE11;
  279: value <= 32'h41858593;
  280: value <= 32'h442295A2;
  281: value <= 32'h449240B2;
  282: value <= 32'h45410612;
  283: value <= 32'hA3990141;
  284: value <= 32'hB7E54641;
  285: value <= 32'h442240B2;
  286: value <= 32'h01414492;
  287: value <= 32'h71398082;
  288: value <= 32'h6985D64E;
  289: value <= 32'hD84ADA26;
  290: value <= 32'h892AD05A;
  291: value <= 32'h41898493;
  292: value <= 32'hD2566B09;
  293: value <= 32'hDE06C86A;
  294: value <= 32'hD452DC22;
  295: value <= 32'hCC62CE5E;
  296: value <= 32'hC66ECA66;
  297: value <= 32'h377994CA;
  298: value <= 32'h99CA4A81;
  299: value <= 32'h0D379B4A;
  300: value <= 32'hA7830100;
  301: value <= 32'hE36340C9;
  302: value <= 32'h153702FA;
  303: value <= 32'h05131A00;
  304: value <= 32'h358DB1C5;
  305: value <= 32'h4109A503;
  306: value <= 32'h153735E1;
  307: value <= 32'h05131A00;
  308: value <= 32'h3D89B185;
  309: value <= 32'h4109A783;
  310: value <= 32'hA0019782;
  311: value <= 32'h1A0017B7;
  312: value <= 32'hB0878513;
  313: value <= 32'h85563581;
  314: value <= 32'h17B73565;
  315: value <= 32'h85131A00;
  316: value <= 32'h3D0DB247;
  317: value <= 32'h0BB740C8;
  318: value <= 32'h4C01E400;
  319: value <= 32'hAA033D51;
  320: value <= 32'hAC830044;
  321: value <= 32'hAD830004;
  322: value <= 32'h9BD20084;
  323: value <= 32'h656344D4;
  324: value <= 32'h0A8500DC;
  325: value <= 32'hBF7104C1;
  326: value <= 32'h920B2403;
  327: value <= 32'h008DF563;
  328: value <= 32'h003D8413;
  329: value <= 32'h86229871;
  330: value <= 32'h01ABFB63;
  331: value <= 32'h856685D2;
  332: value <= 32'h9A222151;
  333: value <= 32'h8DB39CA2;
  334: value <= 32'h0C05408D;
  335: value <= 32'h85CABFC1;
  336: value <= 32'h298D8566;
  337: value <= 32'h85CA8622;
  338: value <= 32'h3E998552;
  339: value <= 32'h882AB7DD;
  340: value <= 32'h4505C57D;
  341: value <= 32'h0EA80863;
  342: value <= 32'h45114889;
  343: value <= 32'h0F181063;
  344: value <= 32'h1A100837;
  345: value <= 32'h04080813;
  346: value <= 32'h450D4891;
  347: value <= 32'h0CB8F863;
  348: value <= 32'hFFF60593;
  349: value <= 32'h81C105C2;
  350: value <= 32'h7FE00893;
  351: value <= 32'hEF634509;
  352: value <= 32'h45BD0AB8;
  353: value <= 32'hEB634505;
  354: value <= 32'h25830AD5;
  355: value <= 32'h05370008;
  356: value <= 32'h8B0D0008;
  357: value <= 32'h20238DC9;
  358: value <= 32'h258300B8;
  359: value <= 32'h05370008;
  360: value <= 32'h157DFFFC;
  361: value <= 32'h0045E593;
  362: value <= 32'h00B82023;
  363: value <= 32'h00082583;
  364: value <= 32'h06120792;
  365: value <= 32'h202399ED;
  366: value <= 32'h258300B8;
  367: value <= 32'h06F20008;
  368: value <= 32'h8DE98E55;
  369: value <= 32'h00B82023;
  370: value <= 32'h00082583;
  371: value <= 32'h20238F4D;
  372: value <= 32'h270300E8;
  373: value <= 32'h8FD90008;
  374: value <= 32'h00F82023;
  375: value <= 32'h00082783;
  376: value <= 32'h00040737;
  377: value <= 32'h00F82023;
  378: value <= 32'h080007B7;
  379: value <= 32'h00082223;
  380: value <= 32'h24238E5D;
  381: value <= 32'h262300C8;
  382: value <= 32'h07930008;
  383: value <= 32'h28230640;
  384: value <= 32'h079300F8;
  385: value <= 32'h2A232690;
  386: value <= 32'h278300F8;
  387: value <= 32'hE7930008;
  388: value <= 32'h20230047;
  389: value <= 32'h278300F8;
  390: value <= 32'h8FD90008;
  391: value <= 32'h00F82023;
  392: value <= 32'h270367C1;
  393: value <= 32'h54630108;
  394: value <= 32'h27830207;
  395: value <= 32'h07370008;
  396: value <= 32'h177DFFF8;
  397: value <= 32'h20238FF9;
  398: value <= 32'h450100F8;
  399: value <= 32'h08378082;
  400: value <= 32'hB71D1A10;
  401: value <= 32'h1A100837;
  402: value <= 32'h02080813;
  403: value <= 32'h17FDBF31;
  404: value <= 32'h4515FBE9;
  405: value <= 32'h71798082;
  406: value <= 32'h47014781;
  407: value <= 32'h06134685;
  408: value <= 32'h45A90280;
  409: value <= 32'hD6064501;
  410: value <= 32'hD226D422;
  411: value <= 32'hCE4ED04A;
  412: value <= 32'h3DF1CC52;
  413: value <= 32'h47014781;
  414: value <= 32'h46514685;
  415: value <= 32'h450545A9;
  416: value <= 32'h470135F9;
  417: value <= 32'h46294685;
  418: value <= 32'h478145A9;
  419: value <= 32'h35C14509;
  420: value <= 32'h1C0107B7;
  421: value <= 32'h4505439C;
  422: value <= 32'h1A1047B7;
  423: value <= 32'h0C47A403;
  424: value <= 32'h3311332D;
  425: value <= 32'h06200793;
  426: value <= 32'h05638805;
  427: value <= 32'h051300F5;
  428: value <= 32'h33010620;
  429: value <= 32'h859365F1;
  430: value <= 32'h45052005;
  431: value <= 32'h1537264D;
  432: value <= 32'h05131A00;
  433: value <= 32'h39B9B2C5;
  434: value <= 32'h1A001537;
  435: value <= 32'hB3850513;
  436: value <= 32'h15373991;
  437: value <= 32'h05131A00;
  438: value <= 32'h31A9B3C5;
  439: value <= 32'h1A001537;
  440: value <= 32'hB4850513;
  441: value <= 32'hC4553181;
  442: value <= 32'h1A001537;
  443: value <= 32'hB6050513;
  444: value <= 32'h25B73915;
  445: value <= 32'h85930026;
  446: value <= 32'h45015A05;
  447: value <= 32'h45812235;
  448: value <= 32'h22ED4501;
  449: value <= 32'h45014581;
  450: value <= 32'h002824A1;
  451: value <= 32'hE4092A91;
  452: value <= 32'h02E00793;
  453: value <= 32'h00F10423;
  454: value <= 32'h000104A3;
  455: value <= 32'hC537C44D;
  456: value <= 32'h67851C07;
  457: value <= 32'h00050413;
  458: value <= 32'h09336489;
  459: value <= 32'h05130094;
  460: value <= 32'h943E0005;
  461: value <= 32'h92F92023;
  462: value <= 32'h90092E23;
  463: value <= 32'h40042223;
  464: value <= 32'h92092223;
  465: value <= 32'h278339C5;
  466: value <= 32'h28039209;
  467: value <= 32'hD73740C4;
  468: value <= 32'h88931C07;
  469: value <= 32'h06B3FFF7;
  470: value <= 32'h071340F0;
  471: value <= 32'h46014207;
  472: value <= 32'h1C000537;
  473: value <= 32'h92848493;
  474: value <= 32'h03061A63;
  475: value <= 32'h97AA6789;
  476: value <= 32'hA0236605;
  477: value <= 32'h061392C7;
  478: value <= 32'h962A5196;
  479: value <= 32'h1A0005B7;
  480: value <= 32'h9007AE23;
  481: value <= 32'h9207A223;
  482: value <= 32'h40060613;
  483: value <= 32'h47E58593;
  484: value <= 32'h15373211;
  485: value <= 32'h05131A00;
  486: value <= 32'hBF99B645;
  487: value <= 32'hFFC72783;
  488: value <= 32'h00F56963;
  489: value <= 32'h95BE430C;
  490: value <= 32'h00B56963;
  491: value <= 32'h07410605;
  492: value <= 32'h05B3BF65;
  493: value <= 32'hFBE30095;
  494: value <= 32'h430CFEB7;
  495: value <= 32'h97C697AE;
  496: value <= 32'h00D7F533;
  497: value <= 32'h345DB7E5;
  498: value <= 32'h1A1047B7;
  499: value <= 32'h0DC7A683;
  500: value <= 32'h05134705;
  501: value <= 32'h88630270;
  502: value <= 32'hA78300E6;
  503: value <= 32'h8B890DC7;
  504: value <= 32'h0513C781;
  505: value <= 32'h31990280;
  506: value <= 32'h1A1047B7;
  507: value <= 32'hDBF84705;
  508: value <= 32'h0007A4B7;
  509: value <= 32'h1A104937;
  510: value <= 32'hEA374985;
  511: value <= 32'h84131C07;
  512: value <= 32'h27831204;
  513: value <= 32'h88630749;
  514: value <= 32'h87B70137;
  515: value <= 32'h87931C00;
  516: value <= 32'h97820807;
  517: value <= 32'h147DA001;
  518: value <= 32'hF46532C1;
  519: value <= 32'hC68A4783;
  520: value <= 32'h0028FFF9;
  521: value <= 32'hBFE13601;
  522: value <= 32'h1A102737;
  523: value <= 32'h47914714;
  524: value <= 32'h00A79533;
  525: value <= 32'hC7148EC9;
  526: value <= 32'h47934714;
  527: value <= 32'h8FF5FFF5;
  528: value <= 32'h431CC71C;
  529: value <= 32'h57B78D5D;
  530: value <= 32'h8793004C;
  531: value <= 32'hD7B3B407;
  532: value <= 32'hC30802B7;
  533: value <= 32'h1C07E737;
  534: value <= 32'h05234501;
  535: value <= 32'h8082C6F7;
  536: value <= 32'h1A102637;
  537: value <= 32'h18864703;
  538: value <= 32'h1C07E6B7;
  539: value <= 32'h18060793;
  540: value <= 32'h04239B3D;
  541: value <= 32'h470318E6;
  542: value <= 32'h9B3D1986;
  543: value <= 32'h18E60C23;
  544: value <= 32'h1A864703;
  545: value <= 32'h04239B3D;
  546: value <= 32'hC6831AE6;
  547: value <= 32'hE737C6A6;
  548: value <= 32'h07131C07;
  549: value <= 32'hC314C287;
  550: value <= 32'h100006B7;
  551: value <= 32'h06B7C354;
  552: value <= 32'h86932007;
  553: value <= 32'hC71409F6;
  554: value <= 32'h704706B7;
  555: value <= 32'hC754068D;
  556: value <= 32'h900006B7;
  557: value <= 32'hCB140685;
  558: value <= 32'h18A62023;
  559: value <= 32'hC3D44691;
  560: value <= 32'h18864683;
  561: value <= 32'h0106E693;
  562: value <= 32'h18D60423;
  563: value <= 32'h4751D398;
  564: value <= 32'h4703D3D8;
  565: value <= 32'h67131A86;
  566: value <= 32'h04230107;
  567: value <= 32'h27371AE6;
  568: value <= 32'h07931A10;
  569: value <= 32'h43DC1807;
  570: value <= 32'h8082FFED;
  571: value <= 32'h003427B7;
  572: value <= 32'h04378793;
  573: value <= 32'h051E953E;
  574: value <= 32'h02854783;
  575: value <= 32'h1C07E737;
  576: value <= 32'hC6A74703;
  577: value <= 32'h04239BBD;
  578: value <= 32'h478302F5;
  579: value <= 32'hE7930285;
  580: value <= 32'h04230407;
  581: value <= 32'hE7B702F5;
  582: value <= 32'h87931C07;
  583: value <= 32'hC398C287;
  584: value <= 32'h10000737;
  585: value <= 32'h07378DD9;
  586: value <= 32'h07132007;
  587: value <= 32'hC7980667;
  588: value <= 32'h90000737;
  589: value <= 32'hD11C0705;
  590: value <= 32'hC7D8C3CC;
  591: value <= 32'hD15C47C1;
  592: value <= 32'h02854783;
  593: value <= 32'h0107E793;
  594: value <= 32'h02F50423;
  595: value <= 32'h80824501;
  596: value <= 32'h003427B7;
  597: value <= 32'h04378793;
  598: value <= 32'h051E953E;
  599: value <= 32'h02854783;
  600: value <= 32'h1C07E737;
  601: value <= 32'hC6A74703;
  602: value <= 32'h04239BBD;
  603: value <= 32'h478302F5;
  604: value <= 32'hE7930285;
  605: value <= 32'h04230407;
  606: value <= 32'hE7B702F5;
  607: value <= 32'h87931C07;
  608: value <= 32'hC398C287;
  609: value <= 32'h10000737;
  610: value <= 32'h07378DD9;
  611: value <= 32'h07132007;
  612: value <= 32'hC7980997;
  613: value <= 32'h90000737;
  614: value <= 32'hD11C0705;
  615: value <= 32'hC7D8C3CC;
  616: value <= 32'hD15C47C1;
  617: value <= 32'h02854783;
  618: value <= 32'h0107E793;
  619: value <= 32'h02F50423;
  620: value <= 32'h80824501;
  621: value <= 32'h1A102837;
  622: value <= 32'h18884703;
  623: value <= 32'h1C07E6B7;
  624: value <= 32'h200708B7;
  625: value <= 32'h04239B3D;
  626: value <= 32'h470318E8;
  627: value <= 32'h03371988;
  628: value <= 32'h0793200F;
  629: value <= 32'h9B3D1808;
  630: value <= 32'h18E80C23;
  631: value <= 32'h1A884703;
  632: value <= 32'h04239B3D;
  633: value <= 32'hC6831AE8;
  634: value <= 32'hE737C6A6;
  635: value <= 32'h07131C07;
  636: value <= 32'hC314C287;
  637: value <= 32'h100006B7;
  638: value <= 32'h8693C354;
  639: value <= 32'hC7140038;
  640: value <= 32'h00855693;
  641: value <= 32'h82C106C2;
  642: value <= 32'h0FF57513;
  643: value <= 32'h0066E6B3;
  644: value <= 32'h01156533;
  645: value <= 32'hCB08C754;
  646: value <= 32'hFFF60693;
  647: value <= 32'h70470537;
  648: value <= 32'hCB548EC9;
  649: value <= 32'h900006B7;
  650: value <= 32'hCF140685;
  651: value <= 32'h18B82023;
  652: value <= 32'h4683C3D0;
  653: value <= 32'hE6931888;
  654: value <= 32'h04230106;
  655: value <= 32'hD39818D8;
  656: value <= 32'hD3D84771;
  657: value <= 32'h1A884703;
  658: value <= 32'h01076713;
  659: value <= 32'h1AE80423;
  660: value <= 32'h1A102737;
  661: value <= 32'h18070793;
  662: value <= 32'hFFED43DC;
  663: value <= 32'h27378082;
  664: value <= 32'h47141A10;
  665: value <= 32'h97B34785;
  666: value <= 32'h8EDD00A7;
  667: value <= 32'h4710C714;
  668: value <= 32'hFFF7C693;
  669: value <= 32'hC7148EF1;
  670: value <= 32'h8FD54314;
  671: value <= 32'h27B7C31C;
  672: value <= 32'h87930034;
  673: value <= 32'h953E0417;
  674: value <= 32'h004C57B7;
  675: value <= 32'hB4078793;
  676: value <= 32'h02B7D7B3;
  677: value <= 32'h07C2051E;
  678: value <= 32'h132383C1;
  679: value <= 32'h515C02F5;
  680: value <= 32'h0067E793;
  681: value <= 32'h515CD15C;
  682: value <= 32'h0107E793;
  683: value <= 32'h515CD15C;
  684: value <= 32'h1007E793;
  685: value <= 32'h515CD15C;
  686: value <= 32'h2007E793;
  687: value <= 32'h4501D15C;
  688: value <= 32'h27B78082;
  689: value <= 32'h87930034;
  690: value <= 32'h953E0417;
  691: value <= 32'h00751793;
  692: value <= 32'h4BD84501;
  693: value <= 32'hCB90EF11;
  694: value <= 32'hC703CBCC;
  695: value <= 32'h67130187;
  696: value <= 32'h8C230107;
  697: value <= 32'h4BD800E7;
  698: value <= 32'h0542E711;
  699: value <= 32'h80828141;
  700: value <= 32'hB7C50505;
  701: value <= 32'hBFC50505;
  702: value <= 32'h4332490A;
  703: value <= 32'h204C4220;
  704: value <= 32'h20504D4A;
  705: value <= 32'h00000000;
  706: value <= 32'h616F4C0A;
  707: value <= 32'h676E6964;
  708: value <= 32'h63655320;
  709: value <= 32'h6E6F6974;
  710: value <= 32'h00000020;
  711: value <= 32'h6D754A0A;
  712: value <= 32'h676E6970;
  713: value <= 32'h206F7420;
  714: value <= 32'h00000000;
  715: value <= 32'h206E614A;
  716: value <= 32'h32203120;
  717: value <= 32'h00323230;
  718: value <= 32'h00002020;
  719: value <= 32'h333A3130;
  720: value <= 32'h38333A31;
  721: value <= 32'h00000000;
  722: value <= 32'h2032410A;
  723: value <= 32'h746F6F42;
  724: value <= 32'h64616F6C;
  725: value <= 32'h42207265;
  726: value <= 32'h73746F6F;
  727: value <= 32'h003D6C65;
  728: value <= 32'h00000031;
  729: value <= 32'h00000030;
  default: value <= 0;
   endcase
  end
endmodule    
